VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM_4k
  CLASS BLOCK ;
  FOREIGN DFFRAM_4k ;
  ORIGIN 0.000 0.000 ;
  SIZE 1694.370 BY 900.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 896.000 26.590 900.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 557.610 896.000 557.890 900.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 610.510 896.000 610.790 900.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 663.870 896.000 664.150 900.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.770 896.000 717.050 900.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 770.130 896.000 770.410 900.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.030 896.000 823.310 900.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.390 896.000 876.670 900.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 896.000 929.570 900.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 982.650 896.000 982.930 900.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1035.550 896.000 1035.830 900.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 896.000 79.490 900.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1088.910 896.000 1089.190 900.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1141.810 896.000 1142.090 900.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 896.000 1195.450 900.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1248.070 896.000 1248.350 900.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1301.430 896.000 1301.710 900.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1354.330 896.000 1354.610 900.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1407.690 896.000 1407.970 900.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1460.590 896.000 1460.870 900.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1513.950 896.000 1514.230 900.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1566.850 896.000 1567.130 900.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 896.000 132.850 900.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1620.210 896.000 1620.490 900.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1673.110 896.000 1673.390 900.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.470 896.000 185.750 900.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 238.830 896.000 239.110 900.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.730 896.000 292.010 900.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.090 896.000 345.370 900.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.990 896.000 398.270 900.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.350 896.000 451.630 900.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.250 896.000 504.530 900.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 823.030 0.000 823.310 4.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1035.550 0.000 1035.830 4.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1088.910 0.000 1089.190 4.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1141.810 0.000 1142.090 4.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1248.070 0.000 1248.350 4.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1301.430 0.000 1301.710 4.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1354.330 0.000 1354.610 4.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1407.690 0.000 1407.970 4.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1460.590 0.000 1460.870 4.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1513.950 0.000 1514.230 4.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.850 0.000 1567.130 4.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.210 0.000 1620.490 4.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.110 0.000 1673.390 4.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.800 4.000 872.400 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1694.180 886.805 ;
      LAYER met1 ;
        RECT 5.520 8.880 1694.180 887.360 ;
      LAYER met2 ;
        RECT 7.000 895.720 26.030 896.000 ;
        RECT 26.870 895.720 78.930 896.000 ;
        RECT 79.770 895.720 132.290 896.000 ;
        RECT 133.130 895.720 185.190 896.000 ;
        RECT 186.030 895.720 238.550 896.000 ;
        RECT 239.390 895.720 291.450 896.000 ;
        RECT 292.290 895.720 344.810 896.000 ;
        RECT 345.650 895.720 397.710 896.000 ;
        RECT 398.550 895.720 451.070 896.000 ;
        RECT 451.910 895.720 503.970 896.000 ;
        RECT 504.810 895.720 557.330 896.000 ;
        RECT 558.170 895.720 610.230 896.000 ;
        RECT 611.070 895.720 663.590 896.000 ;
        RECT 664.430 895.720 716.490 896.000 ;
        RECT 717.330 895.720 769.850 896.000 ;
        RECT 770.690 895.720 822.750 896.000 ;
        RECT 823.590 895.720 876.110 896.000 ;
        RECT 876.950 895.720 929.010 896.000 ;
        RECT 929.850 895.720 982.370 896.000 ;
        RECT 983.210 895.720 1035.270 896.000 ;
        RECT 1036.110 895.720 1088.630 896.000 ;
        RECT 1089.470 895.720 1141.530 896.000 ;
        RECT 1142.370 895.720 1194.890 896.000 ;
        RECT 1195.730 895.720 1247.790 896.000 ;
        RECT 1248.630 895.720 1301.150 896.000 ;
        RECT 1301.990 895.720 1354.050 896.000 ;
        RECT 1354.890 895.720 1407.410 896.000 ;
        RECT 1408.250 895.720 1460.310 896.000 ;
        RECT 1461.150 895.720 1513.670 896.000 ;
        RECT 1514.510 895.720 1566.570 896.000 ;
        RECT 1567.410 895.720 1619.930 896.000 ;
        RECT 1620.770 895.720 1672.830 896.000 ;
        RECT 1673.670 895.720 1691.320 896.000 ;
        RECT 7.000 4.280 1691.320 895.720 ;
        RECT 7.000 4.000 26.030 4.280 ;
        RECT 26.870 4.000 78.930 4.280 ;
        RECT 79.770 4.000 132.290 4.280 ;
        RECT 133.130 4.000 185.190 4.280 ;
        RECT 186.030 4.000 238.550 4.280 ;
        RECT 239.390 4.000 291.450 4.280 ;
        RECT 292.290 4.000 344.810 4.280 ;
        RECT 345.650 4.000 397.710 4.280 ;
        RECT 398.550 4.000 451.070 4.280 ;
        RECT 451.910 4.000 503.970 4.280 ;
        RECT 504.810 4.000 557.330 4.280 ;
        RECT 558.170 4.000 610.230 4.280 ;
        RECT 611.070 4.000 663.590 4.280 ;
        RECT 664.430 4.000 716.490 4.280 ;
        RECT 717.330 4.000 769.850 4.280 ;
        RECT 770.690 4.000 822.750 4.280 ;
        RECT 823.590 4.000 876.110 4.280 ;
        RECT 876.950 4.000 929.010 4.280 ;
        RECT 929.850 4.000 982.370 4.280 ;
        RECT 983.210 4.000 1035.270 4.280 ;
        RECT 1036.110 4.000 1088.630 4.280 ;
        RECT 1089.470 4.000 1141.530 4.280 ;
        RECT 1142.370 4.000 1194.890 4.280 ;
        RECT 1195.730 4.000 1247.790 4.280 ;
        RECT 1248.630 4.000 1301.150 4.280 ;
        RECT 1301.990 4.000 1354.050 4.280 ;
        RECT 1354.890 4.000 1407.410 4.280 ;
        RECT 1408.250 4.000 1460.310 4.280 ;
        RECT 1461.150 4.000 1513.670 4.280 ;
        RECT 1514.510 4.000 1566.570 4.280 ;
        RECT 1567.410 4.000 1619.930 4.280 ;
        RECT 1620.770 4.000 1672.830 4.280 ;
        RECT 1673.670 4.000 1691.320 4.280 ;
      LAYER met3 ;
        RECT 4.000 872.800 1686.295 886.885 ;
        RECT 4.400 871.400 1686.295 872.800 ;
        RECT 4.000 816.360 1686.295 871.400 ;
        RECT 4.400 814.960 1686.295 816.360 ;
        RECT 4.000 759.920 1686.295 814.960 ;
        RECT 4.400 758.520 1686.295 759.920 ;
        RECT 4.000 704.160 1686.295 758.520 ;
        RECT 4.400 702.760 1686.295 704.160 ;
        RECT 4.000 647.720 1686.295 702.760 ;
        RECT 4.400 646.320 1686.295 647.720 ;
        RECT 4.000 591.280 1686.295 646.320 ;
        RECT 4.400 589.880 1686.295 591.280 ;
        RECT 4.000 534.840 1686.295 589.880 ;
        RECT 4.400 533.440 1686.295 534.840 ;
        RECT 4.000 479.080 1686.295 533.440 ;
        RECT 4.400 477.680 1686.295 479.080 ;
        RECT 4.000 422.640 1686.295 477.680 ;
        RECT 4.400 421.240 1686.295 422.640 ;
        RECT 4.000 366.200 1686.295 421.240 ;
        RECT 4.400 364.800 1686.295 366.200 ;
        RECT 4.000 309.760 1686.295 364.800 ;
        RECT 4.400 308.360 1686.295 309.760 ;
        RECT 4.000 254.000 1686.295 308.360 ;
        RECT 4.400 252.600 1686.295 254.000 ;
        RECT 4.000 197.560 1686.295 252.600 ;
        RECT 4.400 196.160 1686.295 197.560 ;
        RECT 4.000 141.120 1686.295 196.160 ;
        RECT 4.400 139.720 1686.295 141.120 ;
        RECT 4.000 84.680 1686.295 139.720 ;
        RECT 4.400 83.280 1686.295 84.680 ;
        RECT 4.000 28.920 1686.295 83.280 ;
        RECT 4.400 27.520 1686.295 28.920 ;
        RECT 4.000 10.715 1686.295 27.520 ;
      LAYER met4 ;
        RECT 29.735 10.640 97.440 886.960 ;
        RECT 99.840 10.640 1675.025 886.960 ;
      LAYER met5 ;
        RECT 1151.500 235.500 1407.020 505.700 ;
  END
END DFFRAM_4k
END LIBRARY

