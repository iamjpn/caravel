VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO register_file_16_1489f923c4dca729178b3e3233458550d8dddf29
  CLASS BLOCK ;
  FOREIGN register_file_16_1489f923c4dca729178b3e3233458550d8dddf29 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1193.470 BY 1204.190 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.970 1200.190 174.250 1204.190 ;
    END
  END clk
  PIN d_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.170 1200.190 1126.450 1204.190 ;
    END
  END d_in[0]
  PIN d_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 1200.190 36.250 1204.190 ;
    END
  END d_in[10]
  PIN d_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 47.640 1193.470 48.240 ;
    END
  END d_in[11]
  PIN d_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END d_in[12]
  PIN d_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END d_in[13]
  PIN d_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1153.770 1200.190 1154.050 1204.190 ;
    END
  END d_in[14]
  PIN d_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END d_in[15]
  PIN d_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END d_in[16]
  PIN d_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 399.880 1193.470 400.480 ;
    END
  END d_in[17]
  PIN d_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END d_in[18]
  PIN d_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1022.760 1193.470 1023.360 ;
    END
  END d_in[19]
  PIN d_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END d_in[1]
  PIN d_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.490 1200.190 823.770 1204.190 ;
    END
  END d_in[20]
  PIN d_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END d_in[21]
  PIN d_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 1200.190 8.650 1204.190 ;
    END
  END d_in[22]
  PIN d_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 590.280 1193.470 590.880 ;
    END
  END d_in[23]
  PIN d_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END d_in[2]
  PIN d_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END d_in[3]
  PIN d_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END d_in[4]
  PIN d_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 658.810 1200.190 659.090 1204.190 ;
    END
  END d_in[5]
  PIN d_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END d_in[6]
  PIN d_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.050 1200.190 357.330 1204.190 ;
    END
  END d_in[7]
  PIN d_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 359.080 1193.470 359.680 ;
    END
  END d_in[8]
  PIN d_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END d_in[9]
  PIN d_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END d_out[0]
  PIN d_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END d_out[100]
  PIN d_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END d_out[101]
  PIN d_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END d_out[102]
  PIN d_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.210 1200.190 631.490 1204.190 ;
    END
  END d_out[103]
  PIN d_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 338.650 1200.190 338.930 1204.190 ;
    END
  END d_out[104]
  PIN d_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 915.490 1200.190 915.770 1204.190 ;
    END
  END d_out[105]
  PIN d_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END d_out[106]
  PIN d_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END d_out[107]
  PIN d_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.530 1200.190 420.810 1204.190 ;
    END
  END d_out[108]
  PIN d_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END d_out[109]
  PIN d_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.530 0.000 1156.810 4.000 ;
    END
  END d_out[10]
  PIN d_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1185.960 1193.470 1186.560 ;
    END
  END d_out[110]
  PIN d_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.690 1200.190 924.970 1204.190 ;
    END
  END d_out[111]
  PIN d_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.930 1200.190 531.210 1204.190 ;
    END
  END d_out[112]
  PIN d_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1052.570 1200.190 1052.850 1204.190 ;
    END
  END d_out[113]
  PIN d_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END d_out[114]
  PIN d_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.370 1200.190 146.650 1204.190 ;
    END
  END d_out[115]
  PIN d_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END d_out[116]
  PIN d_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 792.920 1193.470 793.520 ;
    END
  END d_out[117]
  PIN d_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 375.450 1200.190 375.730 1204.190 ;
    END
  END d_out[118]
  PIN d_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1070.970 1200.190 1071.250 1204.190 ;
    END
  END d_out[119]
  PIN d_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1184.130 0.000 1184.410 4.000 ;
    END
  END d_out[11]
  PIN d_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END d_out[120]
  PIN d_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END d_out[121]
  PIN d_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.330 1200.190 549.610 1204.190 ;
    END
  END d_out[122]
  PIN d_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.880 4.000 1114.480 ;
    END
  END d_out[123]
  PIN d_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1080.170 1200.190 1080.450 1204.190 ;
    END
  END d_out[124]
  PIN d_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END d_out[125]
  PIN d_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END d_out[126]
  PIN d_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 61.240 1193.470 61.840 ;
    END
  END d_out[127]
  PIN d_out[128]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 4.000 ;
    END
  END d_out[128]
  PIN d_out[129]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.130 1200.190 402.410 1204.190 ;
    END
  END d_out[129]
  PIN d_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.450 1200.190 237.730 1204.190 ;
    END
  END d_out[12]
  PIN d_out[130]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 427.080 1193.470 427.680 ;
    END
  END d_out[130]
  PIN d_out[131]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END d_out[131]
  PIN d_out[132]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 841.890 1200.190 842.170 1204.190 ;
    END
  END d_out[132]
  PIN d_out[133]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 890.650 0.000 890.930 4.000 ;
    END
  END d_out[133]
  PIN d_out[134]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1018.530 0.000 1018.810 4.000 ;
    END
  END d_out[134]
  PIN d_out[135]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1104.360 1193.470 1104.960 ;
    END
  END d_out[135]
  PIN d_out[136]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END d_out[136]
  PIN d_out[137]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END d_out[137]
  PIN d_out[138]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END d_out[138]
  PIN d_out[139]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 878.690 1200.190 878.970 1204.190 ;
    END
  END d_out[139]
  PIN d_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.530 1200.190 558.810 1204.190 ;
    END
  END d_out[13]
  PIN d_out[140]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.050 1200.190 311.330 1204.190 ;
    END
  END d_out[140]
  PIN d_out[141]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END d_out[141]
  PIN d_out[142]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 384.650 1200.190 384.930 1204.190 ;
    END
  END d_out[142]
  PIN d_out[143]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END d_out[143]
  PIN d_out[144]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 1200.190 91.450 1204.190 ;
    END
  END d_out[144]
  PIN d_out[145]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END d_out[145]
  PIN d_out[146]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END d_out[146]
  PIN d_out[147]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END d_out[147]
  PIN d_out[148]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END d_out[148]
  PIN d_out[149]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END d_out[149]
  PIN d_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 8.200 1193.470 8.800 ;
    END
  END d_out[14]
  PIN d_out[150]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 952.290 1200.190 952.570 1204.190 ;
    END
  END d_out[150]
  PIN d_out[151]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.330 1200.190 503.610 1204.190 ;
    END
  END d_out[151]
  PIN d_out[152]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 643.320 1193.470 643.920 ;
    END
  END d_out[152]
  PIN d_out[153]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END d_out[153]
  PIN d_out[154]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END d_out[154]
  PIN d_out[155]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END d_out[155]
  PIN d_out[156]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.170 1200.190 183.450 1204.190 ;
    END
  END d_out[156]
  PIN d_out[157]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 918.250 0.000 918.530 4.000 ;
    END
  END d_out[157]
  PIN d_out[158]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END d_out[158]
  PIN d_out[159]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END d_out[159]
  PIN d_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 210.840 1193.470 211.440 ;
    END
  END d_out[15]
  PIN d_out[160]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 851.090 1200.190 851.370 1204.190 ;
    END
  END d_out[160]
  PIN d_out[161]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 4.000 1032.880 ;
    END
  END d_out[161]
  PIN d_out[162]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END d_out[162]
  PIN d_out[163]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END d_out[163]
  PIN d_out[164]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END d_out[164]
  PIN d_out[165]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 265.050 1200.190 265.330 1204.190 ;
    END
  END d_out[165]
  PIN d_out[166]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.330 1200.190 457.610 1204.190 ;
    END
  END d_out[166]
  PIN d_out[167]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END d_out[167]
  PIN d_out[168]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 927.560 1193.470 928.160 ;
    END
  END d_out[168]
  PIN d_out[169]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END d_out[169]
  PIN d_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END d_out[16]
  PIN d_out[170]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.850 1200.190 348.130 1204.190 ;
    END
  END d_out[170]
  PIN d_out[171]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1009.160 1193.470 1009.760 ;
    END
  END d_out[171]
  PIN d_out[172]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 197.240 1193.470 197.840 ;
    END
  END d_out[172]
  PIN d_out[173]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.730 1200.190 476.010 1204.190 ;
    END
  END d_out[173]
  PIN d_out[174]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.280 4.000 964.880 ;
    END
  END d_out[174]
  PIN d_out[175]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1172.170 1200.190 1172.450 1204.190 ;
    END
  END d_out[175]
  PIN d_out[176]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1001.050 0.000 1001.330 4.000 ;
    END
  END d_out[176]
  PIN d_out[177]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.970 1200.190 128.250 1204.190 ;
    END
  END d_out[177]
  PIN d_out[178]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END d_out[178]
  PIN d_out[179]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.050 0.000 909.330 4.000 ;
    END
  END d_out[179]
  PIN d_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END d_out[17]
  PIN d_out[180]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 790.370 0.000 790.650 4.000 ;
    END
  END d_out[180]
  PIN d_out[181]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 888.120 1193.470 888.720 ;
    END
  END d_out[181]
  PIN d_out[182]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 629.720 1193.470 630.320 ;
    END
  END d_out[182]
  PIN d_out[183]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END d_out[183]
  PIN d_out[184]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 209.850 1200.190 210.130 1204.190 ;
    END
  END d_out[184]
  PIN d_out[185]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.080 4.000 1005.680 ;
    END
  END d_out[185]
  PIN d_out[186]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 129.240 1193.470 129.840 ;
    END
  END d_out[186]
  PIN d_out[187]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 535.880 1193.470 536.480 ;
    END
  END d_out[187]
  PIN d_out[188]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1117.960 1193.470 1118.560 ;
    END
  END d_out[188]
  PIN d_out[189]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 301.850 1200.190 302.130 1204.190 ;
    END
  END d_out[189]
  PIN d_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END d_out[18]
  PIN d_out[190]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END d_out[190]
  PIN d_out[191]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END d_out[191]
  PIN d_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END d_out[19]
  PIN d_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 251.640 1193.470 252.240 ;
    END
  END d_out[1]
  PIN d_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 386.280 1193.470 386.880 ;
    END
  END d_out[20]
  PIN d_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END d_out[21]
  PIN d_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 943.090 1200.190 943.370 1204.190 ;
    END
  END d_out[22]
  PIN d_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END d_out[23]
  PIN d_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1181.880 4.000 1182.480 ;
    END
  END d_out[24]
  PIN d_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END d_out[25]
  PIN d_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END d_out[26]
  PIN d_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 292.440 1193.470 293.040 ;
    END
  END d_out[27]
  PIN d_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END d_out[28]
  PIN d_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 567.730 1200.190 568.010 1204.190 ;
    END
  END d_out[29]
  PIN d_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END d_out[2]
  PIN d_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1098.570 1200.190 1098.850 1204.190 ;
    END
  END d_out[30]
  PIN d_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 787.610 1200.190 787.890 1204.190 ;
    END
  END d_out[31]
  PIN d_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 563.080 1193.470 563.680 ;
    END
  END d_out[32]
  PIN d_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 668.010 1200.190 668.290 1204.190 ;
    END
  END d_out[33]
  PIN d_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END d_out[34]
  PIN d_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.930 1200.190 393.210 1204.190 ;
    END
  END d_out[35]
  PIN d_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END d_out[36]
  PIN d_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END d_out[37]
  PIN d_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END d_out[38]
  PIN d_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 765.720 1193.470 766.320 ;
    END
  END d_out[39]
  PIN d_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END d_out[3]
  PIN d_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 752.120 1193.470 752.720 ;
    END
  END d_out[40]
  PIN d_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 440.680 1193.470 441.280 ;
    END
  END d_out[41]
  PIN d_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.770 1200.190 119.050 1204.190 ;
    END
  END d_out[42]
  PIN d_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 995.560 1193.470 996.160 ;
    END
  END d_out[43]
  PIN d_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END d_out[44]
  PIN d_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END d_out[45]
  PIN d_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 494.130 1200.190 494.410 1204.190 ;
    END
  END d_out[46]
  PIN d_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 979.890 1200.190 980.170 1204.190 ;
    END
  END d_out[47]
  PIN d_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 795.890 1200.190 796.170 1204.190 ;
    END
  END d_out[48]
  PIN d_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END d_out[49]
  PIN d_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END d_out[4]
  PIN d_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 981.960 1193.470 982.560 ;
    END
  END d_out[50]
  PIN d_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END d_out[51]
  PIN d_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END d_out[52]
  PIN d_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END d_out[53]
  PIN d_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.530 1200.190 466.810 1204.190 ;
    END
  END d_out[54]
  PIN d_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1089.370 1200.190 1089.650 1204.190 ;
    END
  END d_out[55]
  PIN d_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END d_out[56]
  PIN d_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 686.410 1200.190 686.690 1204.190 ;
    END
  END d_out[57]
  PIN d_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.080 4.000 1073.680 ;
    END
  END d_out[58]
  PIN d_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END d_out[59]
  PIN d_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 711.320 1193.470 711.920 ;
    END
  END d_out[5]
  PIN d_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.610 1200.190 603.890 1204.190 ;
    END
  END d_out[60]
  PIN d_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 741.610 1200.190 741.890 1204.190 ;
    END
  END d_out[61]
  PIN d_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END d_out[62]
  PIN d_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END d_out[63]
  PIN d_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END d_out[64]
  PIN d_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 1200.190 63.850 1204.190 ;
    END
  END d_out[65]
  PIN d_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 833.720 1193.470 834.320 ;
    END
  END d_out[66]
  PIN d_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 941.160 1193.470 941.760 ;
    END
  END d_out[67]
  PIN d_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END d_out[68]
  PIN d_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 901.720 1193.470 902.320 ;
    END
  END d_out[69]
  PIN d_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END d_out[6]
  PIN d_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 156.440 1193.470 157.040 ;
    END
  END d_out[70]
  PIN d_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1100.280 4.000 1100.880 ;
    END
  END d_out[71]
  PIN d_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END d_out[72]
  PIN d_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 714.010 1200.190 714.290 1204.190 ;
    END
  END d_out[73]
  PIN d_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END d_out[74]
  PIN d_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END d_out[75]
  PIN d_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.370 1200.190 997.650 1204.190 ;
    END
  END d_out[76]
  PIN d_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1168.280 4.000 1168.880 ;
    END
  END d_out[77]
  PIN d_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.250 1200.190 320.530 1204.190 ;
    END
  END d_out[78]
  PIN d_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 521.730 1200.190 522.010 1204.190 ;
    END
  END d_out[79]
  PIN d_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.930 1200.190 485.210 1204.190 ;
    END
  END d_out[7]
  PIN d_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 306.040 1193.470 306.640 ;
    END
  END d_out[80]
  PIN d_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 522.280 1193.470 522.880 ;
    END
  END d_out[81]
  PIN d_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END d_out[82]
  PIN d_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1049.960 1193.470 1050.560 ;
    END
  END d_out[83]
  PIN d_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 1200.190 17.850 1204.190 ;
    END
  END d_out[84]
  PIN d_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 684.120 1193.470 684.720 ;
    END
  END d_out[85]
  PIN d_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.080 4.000 1141.680 ;
    END
  END d_out[86]
  PIN d_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.680 4.000 1155.280 ;
    END
  END d_out[87]
  PIN d_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 102.040 1193.470 102.640 ;
    END
  END d_out[88]
  PIN d_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END d_out[89]
  PIN d_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1116.970 1200.190 1117.250 1204.190 ;
    END
  END d_out[8]
  PIN d_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END d_out[90]
  PIN d_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1059.480 4.000 1060.080 ;
    END
  END d_out[91]
  PIN d_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.930 1200.190 439.210 1204.190 ;
    END
  END d_out[92]
  PIN d_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.280 4.000 896.880 ;
    END
  END d_out[93]
  PIN d_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 170.040 1193.470 170.640 ;
    END
  END d_out[94]
  PIN d_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 411.330 1200.190 411.610 1204.190 ;
    END
  END d_out[95]
  PIN d_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END d_out[96]
  PIN d_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END d_out[97]
  PIN d_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END d_out[98]
  PIN d_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1189.650 1200.190 1189.930 1204.190 ;
    END
  END d_out[99]
  PIN d_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 779.320 1193.470 779.920 ;
    END
  END d_out[9]
  PIN dbg_gpr_ack
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 278.840 1193.470 279.440 ;
    END
  END dbg_gpr_ack
  PIN dbg_gpr_addr[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 372.680 1193.470 373.280 ;
    END
  END dbg_gpr_addr[0]
  PIN dbg_gpr_addr[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 887.890 1200.190 888.170 1204.190 ;
    END
  END dbg_gpr_addr[1]
  PIN dbg_gpr_addr[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 142.840 1193.470 143.440 ;
    END
  END dbg_gpr_addr[2]
  PIN dbg_gpr_addr[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 576.680 1193.470 577.280 ;
    END
  END dbg_gpr_addr[3]
  PIN dbg_gpr_addr[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 512.530 1200.190 512.810 1204.190 ;
    END
  END dbg_gpr_addr[4]
  PIN dbg_gpr_addr[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END dbg_gpr_addr[5]
  PIN dbg_gpr_addr[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END dbg_gpr_addr[6]
  PIN dbg_gpr_data[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END dbg_gpr_data[0]
  PIN dbg_gpr_data[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 238.040 1193.470 238.640 ;
    END
  END dbg_gpr_data[10]
  PIN dbg_gpr_data[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END dbg_gpr_data[11]
  PIN dbg_gpr_data[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 115.640 1193.470 116.240 ;
    END
  END dbg_gpr_data[12]
  PIN dbg_gpr_data[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END dbg_gpr_data[13]
  PIN dbg_gpr_data[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 495.080 1193.470 495.680 ;
    END
  END dbg_gpr_data[14]
  PIN dbg_gpr_data[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END dbg_gpr_data[15]
  PIN dbg_gpr_data[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.770 1200.190 165.050 1204.190 ;
    END
  END dbg_gpr_data[16]
  PIN dbg_gpr_data[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 345.480 1193.470 346.080 ;
    END
  END dbg_gpr_data[17]
  PIN dbg_gpr_data[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END dbg_gpr_data[18]
  PIN dbg_gpr_data[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END dbg_gpr_data[19]
  PIN dbg_gpr_data[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 869.490 1200.190 869.770 1204.190 ;
    END
  END dbg_gpr_data[1]
  PIN dbg_gpr_data[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 968.360 1193.470 968.960 ;
    END
  END dbg_gpr_data[20]
  PIN dbg_gpr_data[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END dbg_gpr_data[21]
  PIN dbg_gpr_data[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1119.730 0.000 1120.010 4.000 ;
    END
  END dbg_gpr_data[22]
  PIN dbg_gpr_data[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.290 1200.190 860.570 1204.190 ;
    END
  END dbg_gpr_data[23]
  PIN dbg_gpr_data[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END dbg_gpr_data[24]
  PIN dbg_gpr_data[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END dbg_gpr_data[25]
  PIN dbg_gpr_data[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 413.480 1193.470 414.080 ;
    END
  END dbg_gpr_data[26]
  PIN dbg_gpr_data[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 656.920 1193.470 657.520 ;
    END
  END dbg_gpr_data[27]
  PIN dbg_gpr_data[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END dbg_gpr_data[28]
  PIN dbg_gpr_data[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END dbg_gpr_data[29]
  PIN dbg_gpr_data[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.970 1200.190 1025.250 1204.190 ;
    END
  END dbg_gpr_data[2]
  PIN dbg_gpr_data[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END dbg_gpr_data[30]
  PIN dbg_gpr_data[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END dbg_gpr_data[31]
  PIN dbg_gpr_data[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.880 4.000 978.480 ;
    END
  END dbg_gpr_data[32]
  PIN dbg_gpr_data[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 4.000 ;
    END
  END dbg_gpr_data[33]
  PIN dbg_gpr_data[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END dbg_gpr_data[34]
  PIN dbg_gpr_data[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.250 1200.190 274.530 1204.190 ;
    END
  END dbg_gpr_data[35]
  PIN dbg_gpr_data[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.450 0.000 835.730 4.000 ;
    END
  END dbg_gpr_data[36]
  PIN dbg_gpr_data[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.290 1200.190 814.570 1204.190 ;
    END
  END dbg_gpr_data[37]
  PIN dbg_gpr_data[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 973.450 0.000 973.730 4.000 ;
    END
  END dbg_gpr_data[38]
  PIN dbg_gpr_data[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END dbg_gpr_data[39]
  PIN dbg_gpr_data[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 200.650 1200.190 200.930 1204.190 ;
    END
  END dbg_gpr_data[3]
  PIN dbg_gpr_data[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.130 1200.190 448.410 1204.190 ;
    END
  END dbg_gpr_data[40]
  PIN dbg_gpr_data[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1110.530 0.000 1110.810 4.000 ;
    END
  END dbg_gpr_data[41]
  PIN dbg_gpr_data[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1181.370 1200.190 1181.650 1204.190 ;
    END
  END dbg_gpr_data[42]
  PIN dbg_gpr_data[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1034.170 1200.190 1034.450 1204.190 ;
    END
  END dbg_gpr_data[43]
  PIN dbg_gpr_data[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 594.410 1200.190 594.690 1204.190 ;
    END
  END dbg_gpr_data[44]
  PIN dbg_gpr_data[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.650 1200.190 292.930 1204.190 ;
    END
  END dbg_gpr_data[45]
  PIN dbg_gpr_data[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END dbg_gpr_data[46]
  PIN dbg_gpr_data[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 1200.190 109.850 1204.190 ;
    END
  END dbg_gpr_data[47]
  PIN dbg_gpr_data[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.570 1200.190 155.850 1204.190 ;
    END
  END dbg_gpr_data[48]
  PIN dbg_gpr_data[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END dbg_gpr_data[49]
  PIN dbg_gpr_data[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.880 4.000 1046.480 ;
    END
  END dbg_gpr_data[4]
  PIN dbg_gpr_data[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 954.760 1193.470 955.360 ;
    END
  END dbg_gpr_data[50]
  PIN dbg_gpr_data[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END dbg_gpr_data[51]
  PIN dbg_gpr_data[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 265.240 1193.470 265.840 ;
    END
  END dbg_gpr_data[52]
  PIN dbg_gpr_data[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END dbg_gpr_data[53]
  PIN dbg_gpr_data[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END dbg_gpr_data[54]
  PIN dbg_gpr_data[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 4.000 992.080 ;
    END
  END dbg_gpr_data[55]
  PIN dbg_gpr_data[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END dbg_gpr_data[56]
  PIN dbg_gpr_data[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 454.280 1193.470 454.880 ;
    END
  END dbg_gpr_data[57]
  PIN dbg_gpr_data[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END dbg_gpr_data[58]
  PIN dbg_gpr_data[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1174.930 0.000 1175.210 4.000 ;
    END
  END dbg_gpr_data[59]
  PIN dbg_gpr_data[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 695.610 1200.190 695.890 1204.190 ;
    END
  END dbg_gpr_data[5]
  PIN dbg_gpr_data[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END dbg_gpr_data[60]
  PIN dbg_gpr_data[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.130 1200.190 586.410 1204.190 ;
    END
  END dbg_gpr_data[61]
  PIN dbg_gpr_data[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END dbg_gpr_data[62]
  PIN dbg_gpr_data[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 778.410 1200.190 778.690 1204.190 ;
    END
  END dbg_gpr_data[63]
  PIN dbg_gpr_data[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1145.160 1193.470 1145.760 ;
    END
  END dbg_gpr_data[6]
  PIN dbg_gpr_data[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 255.850 1200.190 256.130 1204.190 ;
    END
  END dbg_gpr_data[7]
  PIN dbg_gpr_data[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 540.130 1200.190 540.410 1204.190 ;
    END
  END dbg_gpr_data[8]
  PIN dbg_gpr_data[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.290 1200.190 906.570 1204.190 ;
    END
  END dbg_gpr_data[9]
  PIN dbg_gpr_req
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 738.520 1193.470 739.120 ;
    END
  END dbg_gpr_req
  PIN log_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1135.370 1200.190 1135.650 1204.190 ;
    END
  END log_out[0]
  PIN log_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END log_out[10]
  PIN log_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1144.570 1200.190 1144.850 1204.190 ;
    END
  END log_out[11]
  PIN log_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.170 1200.190 45.450 1204.190 ;
    END
  END log_out[12]
  PIN log_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 964.250 0.000 964.530 4.000 ;
    END
  END log_out[13]
  PIN log_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 4.000 1194.720 ;
    END
  END log_out[14]
  PIN log_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 616.120 1193.470 616.720 ;
    END
  END log_out[15]
  PIN log_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1036.360 1193.470 1036.960 ;
    END
  END log_out[16]
  PIN log_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 847.320 1193.470 847.920 ;
    END
  END log_out[17]
  PIN log_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END log_out[18]
  PIN log_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 760.010 1200.190 760.290 1204.190 ;
    END
  END log_out[19]
  PIN log_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 74.840 1193.470 75.440 ;
    END
  END log_out[1]
  PIN log_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END log_out[20]
  PIN log_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END log_out[21]
  PIN log_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.370 1200.190 54.650 1204.190 ;
    END
  END log_out[22]
  PIN log_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1127.480 4.000 1128.080 ;
    END
  END log_out[23]
  PIN log_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 897.090 1200.190 897.370 1204.190 ;
    END
  END log_out[24]
  PIN log_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END log_out[25]
  PIN log_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END log_out[26]
  PIN log_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END log_out[27]
  PIN log_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END log_out[28]
  PIN log_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 366.250 1200.190 366.530 1204.190 ;
    END
  END log_out[29]
  PIN log_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END log_out[2]
  PIN log_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END log_out[30]
  PIN log_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END log_out[31]
  PIN log_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 806.520 1193.470 807.120 ;
    END
  END log_out[32]
  PIN log_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 1200.190 73.050 1204.190 ;
    END
  END log_out[33]
  PIN log_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END log_out[34]
  PIN log_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 612.810 1200.190 613.090 1204.190 ;
    END
  END log_out[35]
  PIN log_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END log_out[36]
  PIN log_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 1200.190 137.450 1204.190 ;
    END
  END log_out[37]
  PIN log_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 4.000 951.280 ;
    END
  END log_out[38]
  PIN log_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1172.360 1193.470 1172.960 ;
    END
  END log_out[39]
  PIN log_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END log_out[3]
  PIN log_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END log_out[40]
  PIN log_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.210 1200.190 677.490 1204.190 ;
    END
  END log_out[41]
  PIN log_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 481.480 1193.470 482.080 ;
    END
  END log_out[42]
  PIN log_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END log_out[43]
  PIN log_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1006.570 1200.190 1006.850 1204.190 ;
    END
  END log_out[44]
  PIN log_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END log_out[45]
  PIN log_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 1200.190 27.050 1204.190 ;
    END
  END log_out[46]
  PIN log_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END log_out[47]
  PIN log_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1073.730 0.000 1074.010 4.000 ;
    END
  END log_out[48]
  PIN log_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END log_out[49]
  PIN log_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1101.330 0.000 1101.610 4.000 ;
    END
  END log_out[4]
  PIN log_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 88.440 1193.470 89.040 ;
    END
  END log_out[50]
  PIN log_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END log_out[51]
  PIN log_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END log_out[52]
  PIN log_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.090 1200.190 989.370 1204.190 ;
    END
  END log_out[53]
  PIN log_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 318.280 1193.470 318.880 ;
    END
  END log_out[54]
  PIN log_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 697.720 1193.470 698.320 ;
    END
  END log_out[55]
  PIN log_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 467.880 1193.470 468.480 ;
    END
  END log_out[56]
  PIN log_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END log_out[57]
  PIN log_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 329.450 1200.190 329.730 1204.190 ;
    END
  END log_out[58]
  PIN log_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END log_out[59]
  PIN log_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 183.640 1193.470 184.240 ;
    END
  END log_out[5]
  PIN log_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END log_out[60]
  PIN log_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1063.560 1193.470 1064.160 ;
    END
  END log_out[61]
  PIN log_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END log_out[62]
  PIN log_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END log_out[63]
  PIN log_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 4.000 ;
    END
  END log_out[64]
  PIN log_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.970 1200.190 82.250 1204.190 ;
    END
  END log_out[65]
  PIN log_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 34.040 1193.470 34.640 ;
    END
  END log_out[66]
  PIN log_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.490 1200.190 961.770 1204.190 ;
    END
  END log_out[67]
  PIN log_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1027.730 0.000 1028.010 4.000 ;
    END
  END log_out[68]
  PIN log_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.050 1200.190 219.330 1204.190 ;
    END
  END log_out[69]
  PIN log_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1147.330 0.000 1147.610 4.000 ;
    END
  END log_out[6]
  PIN log_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END log_out[70]
  PIN log_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END log_out[71]
  PIN log_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1131.560 1193.470 1132.160 ;
    END
  END log_out[7]
  PIN log_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1189.470 20.440 1193.470 21.040 ;
    END
  END log_out[8]
  PIN log_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1043.370 1200.190 1043.650 1204.190 ;
    END
  END log_out[9]
  PIN sim_dump
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END sim_dump
  PIN sim_dump_done
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1061.770 1200.190 1062.050 1204.190 ;
    END
  END sim_dump_done
  PIN w_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 508.680 1193.470 509.280 ;
    END
  END w_in[0]
  PIN w_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.010 1200.190 622.290 1204.190 ;
    END
  END w_in[10]
  PIN w_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END w_in[11]
  PIN w_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 283.450 1200.190 283.730 1204.190 ;
    END
  END w_in[12]
  PIN w_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.250 1200.190 228.530 1204.190 ;
    END
  END w_in[13]
  PIN w_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END w_in[14]
  PIN w_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END w_in[15]
  PIN w_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.810 1200.190 705.090 1204.190 ;
    END
  END w_in[16]
  PIN w_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END w_in[17]
  PIN w_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END w_in[18]
  PIN w_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END w_in[19]
  PIN w_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 933.890 1200.190 934.170 1204.190 ;
    END
  END w_in[1]
  PIN w_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1200.190 1108.050 1204.190 ;
    END
  END w_in[20]
  PIN w_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END w_in[21]
  PIN w_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END w_in[22]
  PIN w_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 649.610 1200.190 649.890 1204.190 ;
    END
  END w_in[23]
  PIN w_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END w_in[24]
  PIN w_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 832.690 1200.190 832.970 1204.190 ;
    END
  END w_in[25]
  PIN w_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END w_in[26]
  PIN w_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1086.680 4.000 1087.280 ;
    END
  END w_in[27]
  PIN w_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.930 0.000 1083.210 4.000 ;
    END
  END w_in[28]
  PIN w_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END w_in[29]
  PIN w_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END w_in[2]
  PIN w_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END w_in[30]
  PIN w_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END w_in[31]
  PIN w_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END w_in[32]
  PIN w_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1077.160 1193.470 1077.760 ;
    END
  END w_in[33]
  PIN w_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END w_in[34]
  PIN w_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END w_in[35]
  PIN w_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END w_in[36]
  PIN w_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.330 0.000 1055.610 4.000 ;
    END
  END w_in[37]
  PIN w_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 724.920 1193.470 725.520 ;
    END
  END w_in[38]
  PIN w_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END w_in[39]
  PIN w_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 549.480 1193.470 550.080 ;
    END
  END w_in[3]
  PIN w_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 429.730 1200.190 430.010 1204.190 ;
    END
  END w_in[40]
  PIN w_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 860.920 1193.470 861.520 ;
    END
  END w_in[41]
  PIN w_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END w_in[42]
  PIN w_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 874.520 1193.470 875.120 ;
    END
  END w_in[43]
  PIN w_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 1200.190 100.650 1204.190 ;
    END
  END w_in[44]
  PIN w_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 224.440 1193.470 225.040 ;
    END
  END w_in[45]
  PIN w_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1090.760 1193.470 1091.360 ;
    END
  END w_in[46]
  PIN w_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 1158.760 1193.470 1159.360 ;
    END
  END w_in[47]
  PIN w_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 723.210 1200.190 723.490 1204.190 ;
    END
  END w_in[48]
  PIN w_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END w_in[49]
  PIN w_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1015.770 1200.190 1016.050 1204.190 ;
    END
  END w_in[4]
  PIN w_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.970 1200.190 1163.250 1204.190 ;
    END
  END w_in[50]
  PIN w_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END w_in[51]
  PIN w_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 970.690 1200.190 970.970 1204.190 ;
    END
  END w_in[52]
  PIN w_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END w_in[53]
  PIN w_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 913.960 1193.470 914.560 ;
    END
  END w_in[54]
  PIN w_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.650 1200.190 246.930 1204.190 ;
    END
  END w_in[55]
  PIN w_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.210 1200.190 769.490 1204.190 ;
    END
  END w_in[56]
  PIN w_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END w_in[57]
  PIN w_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END w_in[58]
  PIN w_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 670.520 1193.470 671.120 ;
    END
  END w_in[59]
  PIN w_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END w_in[5]
  PIN w_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 820.120 1193.470 820.720 ;
    END
  END w_in[60]
  PIN w_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 853.850 0.000 854.130 4.000 ;
    END
  END w_in[61]
  PIN w_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END w_in[62]
  PIN w_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END w_in[63]
  PIN w_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 331.880 1193.470 332.480 ;
    END
  END w_in[64]
  PIN w_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1189.470 603.880 1193.470 604.480 ;
    END
  END w_in[65]
  PIN w_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END w_in[66]
  PIN w_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END w_in[67]
  PIN w_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.090 1200.190 805.370 1204.190 ;
    END
  END w_in[68]
  PIN w_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END w_in[69]
  PIN w_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 725.970 0.000 726.250 4.000 ;
    END
  END w_in[6]
  PIN w_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 750.810 1200.190 751.090 1204.190 ;
    END
  END w_in[70]
  PIN w_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 576.930 1200.190 577.210 1204.190 ;
    END
  END w_in[71]
  PIN w_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.450 1200.190 191.730 1204.190 ;
    END
  END w_in[7]
  PIN w_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 732.410 1200.190 732.690 1204.190 ;
    END
  END w_in[8]
  PIN w_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 640.410 1200.190 640.690 1204.190 ;
    END
  END w_in[9]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1191.600 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1191.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1187.720 1191.445 ;
      LAYER met1 ;
        RECT 2.830 4.460 1187.720 1193.700 ;
      LAYER met2 ;
        RECT 2.860 1199.910 8.090 1200.190 ;
        RECT 8.930 1199.910 17.290 1200.190 ;
        RECT 18.130 1199.910 26.490 1200.190 ;
        RECT 27.330 1199.910 35.690 1200.190 ;
        RECT 36.530 1199.910 44.890 1200.190 ;
        RECT 45.730 1199.910 54.090 1200.190 ;
        RECT 54.930 1199.910 63.290 1200.190 ;
        RECT 64.130 1199.910 72.490 1200.190 ;
        RECT 73.330 1199.910 81.690 1200.190 ;
        RECT 82.530 1199.910 90.890 1200.190 ;
        RECT 91.730 1199.910 100.090 1200.190 ;
        RECT 100.930 1199.910 109.290 1200.190 ;
        RECT 110.130 1199.910 118.490 1200.190 ;
        RECT 119.330 1199.910 127.690 1200.190 ;
        RECT 128.530 1199.910 136.890 1200.190 ;
        RECT 137.730 1199.910 146.090 1200.190 ;
        RECT 146.930 1199.910 155.290 1200.190 ;
        RECT 156.130 1199.910 164.490 1200.190 ;
        RECT 165.330 1199.910 173.690 1200.190 ;
        RECT 174.530 1199.910 182.890 1200.190 ;
        RECT 183.730 1199.910 191.170 1200.190 ;
        RECT 192.010 1199.910 200.370 1200.190 ;
        RECT 201.210 1199.910 209.570 1200.190 ;
        RECT 210.410 1199.910 218.770 1200.190 ;
        RECT 219.610 1199.910 227.970 1200.190 ;
        RECT 228.810 1199.910 237.170 1200.190 ;
        RECT 238.010 1199.910 246.370 1200.190 ;
        RECT 247.210 1199.910 255.570 1200.190 ;
        RECT 256.410 1199.910 264.770 1200.190 ;
        RECT 265.610 1199.910 273.970 1200.190 ;
        RECT 274.810 1199.910 283.170 1200.190 ;
        RECT 284.010 1199.910 292.370 1200.190 ;
        RECT 293.210 1199.910 301.570 1200.190 ;
        RECT 302.410 1199.910 310.770 1200.190 ;
        RECT 311.610 1199.910 319.970 1200.190 ;
        RECT 320.810 1199.910 329.170 1200.190 ;
        RECT 330.010 1199.910 338.370 1200.190 ;
        RECT 339.210 1199.910 347.570 1200.190 ;
        RECT 348.410 1199.910 356.770 1200.190 ;
        RECT 357.610 1199.910 365.970 1200.190 ;
        RECT 366.810 1199.910 375.170 1200.190 ;
        RECT 376.010 1199.910 384.370 1200.190 ;
        RECT 385.210 1199.910 392.650 1200.190 ;
        RECT 393.490 1199.910 401.850 1200.190 ;
        RECT 402.690 1199.910 411.050 1200.190 ;
        RECT 411.890 1199.910 420.250 1200.190 ;
        RECT 421.090 1199.910 429.450 1200.190 ;
        RECT 430.290 1199.910 438.650 1200.190 ;
        RECT 439.490 1199.910 447.850 1200.190 ;
        RECT 448.690 1199.910 457.050 1200.190 ;
        RECT 457.890 1199.910 466.250 1200.190 ;
        RECT 467.090 1199.910 475.450 1200.190 ;
        RECT 476.290 1199.910 484.650 1200.190 ;
        RECT 485.490 1199.910 493.850 1200.190 ;
        RECT 494.690 1199.910 503.050 1200.190 ;
        RECT 503.890 1199.910 512.250 1200.190 ;
        RECT 513.090 1199.910 521.450 1200.190 ;
        RECT 522.290 1199.910 530.650 1200.190 ;
        RECT 531.490 1199.910 539.850 1200.190 ;
        RECT 540.690 1199.910 549.050 1200.190 ;
        RECT 549.890 1199.910 558.250 1200.190 ;
        RECT 559.090 1199.910 567.450 1200.190 ;
        RECT 568.290 1199.910 576.650 1200.190 ;
        RECT 577.490 1199.910 585.850 1200.190 ;
        RECT 586.690 1199.910 594.130 1200.190 ;
        RECT 594.970 1199.910 603.330 1200.190 ;
        RECT 604.170 1199.910 612.530 1200.190 ;
        RECT 613.370 1199.910 621.730 1200.190 ;
        RECT 622.570 1199.910 630.930 1200.190 ;
        RECT 631.770 1199.910 640.130 1200.190 ;
        RECT 640.970 1199.910 649.330 1200.190 ;
        RECT 650.170 1199.910 658.530 1200.190 ;
        RECT 659.370 1199.910 667.730 1200.190 ;
        RECT 668.570 1199.910 676.930 1200.190 ;
        RECT 677.770 1199.910 686.130 1200.190 ;
        RECT 686.970 1199.910 695.330 1200.190 ;
        RECT 696.170 1199.910 704.530 1200.190 ;
        RECT 705.370 1199.910 713.730 1200.190 ;
        RECT 714.570 1199.910 722.930 1200.190 ;
        RECT 723.770 1199.910 732.130 1200.190 ;
        RECT 732.970 1199.910 741.330 1200.190 ;
        RECT 742.170 1199.910 750.530 1200.190 ;
        RECT 751.370 1199.910 759.730 1200.190 ;
        RECT 760.570 1199.910 768.930 1200.190 ;
        RECT 769.770 1199.910 778.130 1200.190 ;
        RECT 778.970 1199.910 787.330 1200.190 ;
        RECT 788.170 1199.910 795.610 1200.190 ;
        RECT 796.450 1199.910 804.810 1200.190 ;
        RECT 805.650 1199.910 814.010 1200.190 ;
        RECT 814.850 1199.910 823.210 1200.190 ;
        RECT 824.050 1199.910 832.410 1200.190 ;
        RECT 833.250 1199.910 841.610 1200.190 ;
        RECT 842.450 1199.910 850.810 1200.190 ;
        RECT 851.650 1199.910 860.010 1200.190 ;
        RECT 860.850 1199.910 869.210 1200.190 ;
        RECT 870.050 1199.910 878.410 1200.190 ;
        RECT 879.250 1199.910 887.610 1200.190 ;
        RECT 888.450 1199.910 896.810 1200.190 ;
        RECT 897.650 1199.910 906.010 1200.190 ;
        RECT 906.850 1199.910 915.210 1200.190 ;
        RECT 916.050 1199.910 924.410 1200.190 ;
        RECT 925.250 1199.910 933.610 1200.190 ;
        RECT 934.450 1199.910 942.810 1200.190 ;
        RECT 943.650 1199.910 952.010 1200.190 ;
        RECT 952.850 1199.910 961.210 1200.190 ;
        RECT 962.050 1199.910 970.410 1200.190 ;
        RECT 971.250 1199.910 979.610 1200.190 ;
        RECT 980.450 1199.910 988.810 1200.190 ;
        RECT 989.650 1199.910 997.090 1200.190 ;
        RECT 997.930 1199.910 1006.290 1200.190 ;
        RECT 1007.130 1199.910 1015.490 1200.190 ;
        RECT 1016.330 1199.910 1024.690 1200.190 ;
        RECT 1025.530 1199.910 1033.890 1200.190 ;
        RECT 1034.730 1199.910 1043.090 1200.190 ;
        RECT 1043.930 1199.910 1052.290 1200.190 ;
        RECT 1053.130 1199.910 1061.490 1200.190 ;
        RECT 1062.330 1199.910 1070.690 1200.190 ;
        RECT 1071.530 1199.910 1079.890 1200.190 ;
        RECT 1080.730 1199.910 1089.090 1200.190 ;
        RECT 1089.930 1199.910 1098.290 1200.190 ;
        RECT 1099.130 1199.910 1107.490 1200.190 ;
        RECT 1108.330 1199.910 1116.690 1200.190 ;
        RECT 1117.530 1199.910 1125.890 1200.190 ;
        RECT 1126.730 1199.910 1135.090 1200.190 ;
        RECT 1135.930 1199.910 1144.290 1200.190 ;
        RECT 1145.130 1199.910 1153.490 1200.190 ;
        RECT 1154.330 1199.910 1162.690 1200.190 ;
        RECT 1163.530 1199.910 1171.890 1200.190 ;
        RECT 1172.730 1199.910 1181.090 1200.190 ;
        RECT 1181.930 1199.910 1189.370 1200.190 ;
        RECT 2.860 4.280 1189.930 1199.910 ;
        RECT 3.410 4.000 10.850 4.280 ;
        RECT 11.690 4.000 20.050 4.280 ;
        RECT 20.890 4.000 29.250 4.280 ;
        RECT 30.090 4.000 38.450 4.280 ;
        RECT 39.290 4.000 47.650 4.280 ;
        RECT 48.490 4.000 56.850 4.280 ;
        RECT 57.690 4.000 66.050 4.280 ;
        RECT 66.890 4.000 75.250 4.280 ;
        RECT 76.090 4.000 84.450 4.280 ;
        RECT 85.290 4.000 93.650 4.280 ;
        RECT 94.490 4.000 102.850 4.280 ;
        RECT 103.690 4.000 112.050 4.280 ;
        RECT 112.890 4.000 121.250 4.280 ;
        RECT 122.090 4.000 130.450 4.280 ;
        RECT 131.290 4.000 139.650 4.280 ;
        RECT 140.490 4.000 148.850 4.280 ;
        RECT 149.690 4.000 158.050 4.280 ;
        RECT 158.890 4.000 167.250 4.280 ;
        RECT 168.090 4.000 176.450 4.280 ;
        RECT 177.290 4.000 185.650 4.280 ;
        RECT 186.490 4.000 194.850 4.280 ;
        RECT 195.690 4.000 203.130 4.280 ;
        RECT 203.970 4.000 212.330 4.280 ;
        RECT 213.170 4.000 221.530 4.280 ;
        RECT 222.370 4.000 230.730 4.280 ;
        RECT 231.570 4.000 239.930 4.280 ;
        RECT 240.770 4.000 249.130 4.280 ;
        RECT 249.970 4.000 258.330 4.280 ;
        RECT 259.170 4.000 267.530 4.280 ;
        RECT 268.370 4.000 276.730 4.280 ;
        RECT 277.570 4.000 285.930 4.280 ;
        RECT 286.770 4.000 295.130 4.280 ;
        RECT 295.970 4.000 304.330 4.280 ;
        RECT 305.170 4.000 313.530 4.280 ;
        RECT 314.370 4.000 322.730 4.280 ;
        RECT 323.570 4.000 331.930 4.280 ;
        RECT 332.770 4.000 341.130 4.280 ;
        RECT 341.970 4.000 350.330 4.280 ;
        RECT 351.170 4.000 359.530 4.280 ;
        RECT 360.370 4.000 368.730 4.280 ;
        RECT 369.570 4.000 377.930 4.280 ;
        RECT 378.770 4.000 387.130 4.280 ;
        RECT 387.970 4.000 396.330 4.280 ;
        RECT 397.170 4.000 404.610 4.280 ;
        RECT 405.450 4.000 413.810 4.280 ;
        RECT 414.650 4.000 423.010 4.280 ;
        RECT 423.850 4.000 432.210 4.280 ;
        RECT 433.050 4.000 441.410 4.280 ;
        RECT 442.250 4.000 450.610 4.280 ;
        RECT 451.450 4.000 459.810 4.280 ;
        RECT 460.650 4.000 469.010 4.280 ;
        RECT 469.850 4.000 478.210 4.280 ;
        RECT 479.050 4.000 487.410 4.280 ;
        RECT 488.250 4.000 496.610 4.280 ;
        RECT 497.450 4.000 505.810 4.280 ;
        RECT 506.650 4.000 515.010 4.280 ;
        RECT 515.850 4.000 524.210 4.280 ;
        RECT 525.050 4.000 533.410 4.280 ;
        RECT 534.250 4.000 542.610 4.280 ;
        RECT 543.450 4.000 551.810 4.280 ;
        RECT 552.650 4.000 561.010 4.280 ;
        RECT 561.850 4.000 570.210 4.280 ;
        RECT 571.050 4.000 579.410 4.280 ;
        RECT 580.250 4.000 588.610 4.280 ;
        RECT 589.450 4.000 597.810 4.280 ;
        RECT 598.650 4.000 606.090 4.280 ;
        RECT 606.930 4.000 615.290 4.280 ;
        RECT 616.130 4.000 624.490 4.280 ;
        RECT 625.330 4.000 633.690 4.280 ;
        RECT 634.530 4.000 642.890 4.280 ;
        RECT 643.730 4.000 652.090 4.280 ;
        RECT 652.930 4.000 661.290 4.280 ;
        RECT 662.130 4.000 670.490 4.280 ;
        RECT 671.330 4.000 679.690 4.280 ;
        RECT 680.530 4.000 688.890 4.280 ;
        RECT 689.730 4.000 698.090 4.280 ;
        RECT 698.930 4.000 707.290 4.280 ;
        RECT 708.130 4.000 716.490 4.280 ;
        RECT 717.330 4.000 725.690 4.280 ;
        RECT 726.530 4.000 734.890 4.280 ;
        RECT 735.730 4.000 744.090 4.280 ;
        RECT 744.930 4.000 753.290 4.280 ;
        RECT 754.130 4.000 762.490 4.280 ;
        RECT 763.330 4.000 771.690 4.280 ;
        RECT 772.530 4.000 780.890 4.280 ;
        RECT 781.730 4.000 790.090 4.280 ;
        RECT 790.930 4.000 799.290 4.280 ;
        RECT 800.130 4.000 807.570 4.280 ;
        RECT 808.410 4.000 816.770 4.280 ;
        RECT 817.610 4.000 825.970 4.280 ;
        RECT 826.810 4.000 835.170 4.280 ;
        RECT 836.010 4.000 844.370 4.280 ;
        RECT 845.210 4.000 853.570 4.280 ;
        RECT 854.410 4.000 862.770 4.280 ;
        RECT 863.610 4.000 871.970 4.280 ;
        RECT 872.810 4.000 881.170 4.280 ;
        RECT 882.010 4.000 890.370 4.280 ;
        RECT 891.210 4.000 899.570 4.280 ;
        RECT 900.410 4.000 908.770 4.280 ;
        RECT 909.610 4.000 917.970 4.280 ;
        RECT 918.810 4.000 927.170 4.280 ;
        RECT 928.010 4.000 936.370 4.280 ;
        RECT 937.210 4.000 945.570 4.280 ;
        RECT 946.410 4.000 954.770 4.280 ;
        RECT 955.610 4.000 963.970 4.280 ;
        RECT 964.810 4.000 973.170 4.280 ;
        RECT 974.010 4.000 982.370 4.280 ;
        RECT 983.210 4.000 991.570 4.280 ;
        RECT 992.410 4.000 1000.770 4.280 ;
        RECT 1001.610 4.000 1009.050 4.280 ;
        RECT 1009.890 4.000 1018.250 4.280 ;
        RECT 1019.090 4.000 1027.450 4.280 ;
        RECT 1028.290 4.000 1036.650 4.280 ;
        RECT 1037.490 4.000 1045.850 4.280 ;
        RECT 1046.690 4.000 1055.050 4.280 ;
        RECT 1055.890 4.000 1064.250 4.280 ;
        RECT 1065.090 4.000 1073.450 4.280 ;
        RECT 1074.290 4.000 1082.650 4.280 ;
        RECT 1083.490 4.000 1091.850 4.280 ;
        RECT 1092.690 4.000 1101.050 4.280 ;
        RECT 1101.890 4.000 1110.250 4.280 ;
        RECT 1111.090 4.000 1119.450 4.280 ;
        RECT 1120.290 4.000 1128.650 4.280 ;
        RECT 1129.490 4.000 1137.850 4.280 ;
        RECT 1138.690 4.000 1147.050 4.280 ;
        RECT 1147.890 4.000 1156.250 4.280 ;
        RECT 1157.090 4.000 1165.450 4.280 ;
        RECT 1166.290 4.000 1174.650 4.280 ;
        RECT 1175.490 4.000 1183.850 4.280 ;
        RECT 1184.690 4.000 1189.930 4.280 ;
      LAYER met3 ;
        RECT 4.400 1193.720 1189.955 1194.585 ;
        RECT 3.990 1186.960 1189.955 1193.720 ;
        RECT 3.990 1185.560 1189.070 1186.960 ;
        RECT 3.990 1182.880 1189.955 1185.560 ;
        RECT 4.400 1181.480 1189.955 1182.880 ;
        RECT 3.990 1173.360 1189.955 1181.480 ;
        RECT 3.990 1171.960 1189.070 1173.360 ;
        RECT 3.990 1169.280 1189.955 1171.960 ;
        RECT 4.400 1167.880 1189.955 1169.280 ;
        RECT 3.990 1159.760 1189.955 1167.880 ;
        RECT 3.990 1158.360 1189.070 1159.760 ;
        RECT 3.990 1155.680 1189.955 1158.360 ;
        RECT 4.400 1154.280 1189.955 1155.680 ;
        RECT 3.990 1146.160 1189.955 1154.280 ;
        RECT 3.990 1144.760 1189.070 1146.160 ;
        RECT 3.990 1142.080 1189.955 1144.760 ;
        RECT 4.400 1140.680 1189.955 1142.080 ;
        RECT 3.990 1132.560 1189.955 1140.680 ;
        RECT 3.990 1131.160 1189.070 1132.560 ;
        RECT 3.990 1128.480 1189.955 1131.160 ;
        RECT 4.400 1127.080 1189.955 1128.480 ;
        RECT 3.990 1118.960 1189.955 1127.080 ;
        RECT 3.990 1117.560 1189.070 1118.960 ;
        RECT 3.990 1114.880 1189.955 1117.560 ;
        RECT 4.400 1113.480 1189.955 1114.880 ;
        RECT 3.990 1105.360 1189.955 1113.480 ;
        RECT 3.990 1103.960 1189.070 1105.360 ;
        RECT 3.990 1101.280 1189.955 1103.960 ;
        RECT 4.400 1099.880 1189.955 1101.280 ;
        RECT 3.990 1091.760 1189.955 1099.880 ;
        RECT 3.990 1090.360 1189.070 1091.760 ;
        RECT 3.990 1087.680 1189.955 1090.360 ;
        RECT 4.400 1086.280 1189.955 1087.680 ;
        RECT 3.990 1078.160 1189.955 1086.280 ;
        RECT 3.990 1076.760 1189.070 1078.160 ;
        RECT 3.990 1074.080 1189.955 1076.760 ;
        RECT 4.400 1072.680 1189.955 1074.080 ;
        RECT 3.990 1064.560 1189.955 1072.680 ;
        RECT 3.990 1063.160 1189.070 1064.560 ;
        RECT 3.990 1060.480 1189.955 1063.160 ;
        RECT 4.400 1059.080 1189.955 1060.480 ;
        RECT 3.990 1050.960 1189.955 1059.080 ;
        RECT 3.990 1049.560 1189.070 1050.960 ;
        RECT 3.990 1046.880 1189.955 1049.560 ;
        RECT 4.400 1045.480 1189.955 1046.880 ;
        RECT 3.990 1037.360 1189.955 1045.480 ;
        RECT 3.990 1035.960 1189.070 1037.360 ;
        RECT 3.990 1033.280 1189.955 1035.960 ;
        RECT 4.400 1031.880 1189.955 1033.280 ;
        RECT 3.990 1023.760 1189.955 1031.880 ;
        RECT 3.990 1022.360 1189.070 1023.760 ;
        RECT 3.990 1019.680 1189.955 1022.360 ;
        RECT 4.400 1018.280 1189.955 1019.680 ;
        RECT 3.990 1010.160 1189.955 1018.280 ;
        RECT 3.990 1008.760 1189.070 1010.160 ;
        RECT 3.990 1006.080 1189.955 1008.760 ;
        RECT 4.400 1004.680 1189.955 1006.080 ;
        RECT 3.990 996.560 1189.955 1004.680 ;
        RECT 3.990 995.160 1189.070 996.560 ;
        RECT 3.990 992.480 1189.955 995.160 ;
        RECT 4.400 991.080 1189.955 992.480 ;
        RECT 3.990 982.960 1189.955 991.080 ;
        RECT 3.990 981.560 1189.070 982.960 ;
        RECT 3.990 978.880 1189.955 981.560 ;
        RECT 4.400 977.480 1189.955 978.880 ;
        RECT 3.990 969.360 1189.955 977.480 ;
        RECT 3.990 967.960 1189.070 969.360 ;
        RECT 3.990 965.280 1189.955 967.960 ;
        RECT 4.400 963.880 1189.955 965.280 ;
        RECT 3.990 955.760 1189.955 963.880 ;
        RECT 3.990 954.360 1189.070 955.760 ;
        RECT 3.990 951.680 1189.955 954.360 ;
        RECT 4.400 950.280 1189.955 951.680 ;
        RECT 3.990 942.160 1189.955 950.280 ;
        RECT 3.990 940.760 1189.070 942.160 ;
        RECT 3.990 938.080 1189.955 940.760 ;
        RECT 4.400 936.680 1189.955 938.080 ;
        RECT 3.990 928.560 1189.955 936.680 ;
        RECT 3.990 927.160 1189.070 928.560 ;
        RECT 3.990 924.480 1189.955 927.160 ;
        RECT 4.400 923.080 1189.955 924.480 ;
        RECT 3.990 914.960 1189.955 923.080 ;
        RECT 3.990 913.560 1189.070 914.960 ;
        RECT 3.990 910.880 1189.955 913.560 ;
        RECT 4.400 909.480 1189.955 910.880 ;
        RECT 3.990 902.720 1189.955 909.480 ;
        RECT 3.990 901.320 1189.070 902.720 ;
        RECT 3.990 897.280 1189.955 901.320 ;
        RECT 4.400 895.880 1189.955 897.280 ;
        RECT 3.990 889.120 1189.955 895.880 ;
        RECT 3.990 887.720 1189.070 889.120 ;
        RECT 3.990 885.040 1189.955 887.720 ;
        RECT 4.400 883.640 1189.955 885.040 ;
        RECT 3.990 875.520 1189.955 883.640 ;
        RECT 3.990 874.120 1189.070 875.520 ;
        RECT 3.990 871.440 1189.955 874.120 ;
        RECT 4.400 870.040 1189.955 871.440 ;
        RECT 3.990 861.920 1189.955 870.040 ;
        RECT 3.990 860.520 1189.070 861.920 ;
        RECT 3.990 857.840 1189.955 860.520 ;
        RECT 4.400 856.440 1189.955 857.840 ;
        RECT 3.990 848.320 1189.955 856.440 ;
        RECT 3.990 846.920 1189.070 848.320 ;
        RECT 3.990 844.240 1189.955 846.920 ;
        RECT 4.400 842.840 1189.955 844.240 ;
        RECT 3.990 834.720 1189.955 842.840 ;
        RECT 3.990 833.320 1189.070 834.720 ;
        RECT 3.990 830.640 1189.955 833.320 ;
        RECT 4.400 829.240 1189.955 830.640 ;
        RECT 3.990 821.120 1189.955 829.240 ;
        RECT 3.990 819.720 1189.070 821.120 ;
        RECT 3.990 817.040 1189.955 819.720 ;
        RECT 4.400 815.640 1189.955 817.040 ;
        RECT 3.990 807.520 1189.955 815.640 ;
        RECT 3.990 806.120 1189.070 807.520 ;
        RECT 3.990 803.440 1189.955 806.120 ;
        RECT 4.400 802.040 1189.955 803.440 ;
        RECT 3.990 793.920 1189.955 802.040 ;
        RECT 3.990 792.520 1189.070 793.920 ;
        RECT 3.990 789.840 1189.955 792.520 ;
        RECT 4.400 788.440 1189.955 789.840 ;
        RECT 3.990 780.320 1189.955 788.440 ;
        RECT 3.990 778.920 1189.070 780.320 ;
        RECT 3.990 776.240 1189.955 778.920 ;
        RECT 4.400 774.840 1189.955 776.240 ;
        RECT 3.990 766.720 1189.955 774.840 ;
        RECT 3.990 765.320 1189.070 766.720 ;
        RECT 3.990 762.640 1189.955 765.320 ;
        RECT 4.400 761.240 1189.955 762.640 ;
        RECT 3.990 753.120 1189.955 761.240 ;
        RECT 3.990 751.720 1189.070 753.120 ;
        RECT 3.990 749.040 1189.955 751.720 ;
        RECT 4.400 747.640 1189.955 749.040 ;
        RECT 3.990 739.520 1189.955 747.640 ;
        RECT 3.990 738.120 1189.070 739.520 ;
        RECT 3.990 735.440 1189.955 738.120 ;
        RECT 4.400 734.040 1189.955 735.440 ;
        RECT 3.990 725.920 1189.955 734.040 ;
        RECT 3.990 724.520 1189.070 725.920 ;
        RECT 3.990 721.840 1189.955 724.520 ;
        RECT 4.400 720.440 1189.955 721.840 ;
        RECT 3.990 712.320 1189.955 720.440 ;
        RECT 3.990 710.920 1189.070 712.320 ;
        RECT 3.990 708.240 1189.955 710.920 ;
        RECT 4.400 706.840 1189.955 708.240 ;
        RECT 3.990 698.720 1189.955 706.840 ;
        RECT 3.990 697.320 1189.070 698.720 ;
        RECT 3.990 694.640 1189.955 697.320 ;
        RECT 4.400 693.240 1189.955 694.640 ;
        RECT 3.990 685.120 1189.955 693.240 ;
        RECT 3.990 683.720 1189.070 685.120 ;
        RECT 3.990 681.040 1189.955 683.720 ;
        RECT 4.400 679.640 1189.955 681.040 ;
        RECT 3.990 671.520 1189.955 679.640 ;
        RECT 3.990 670.120 1189.070 671.520 ;
        RECT 3.990 667.440 1189.955 670.120 ;
        RECT 4.400 666.040 1189.955 667.440 ;
        RECT 3.990 657.920 1189.955 666.040 ;
        RECT 3.990 656.520 1189.070 657.920 ;
        RECT 3.990 653.840 1189.955 656.520 ;
        RECT 4.400 652.440 1189.955 653.840 ;
        RECT 3.990 644.320 1189.955 652.440 ;
        RECT 3.990 642.920 1189.070 644.320 ;
        RECT 3.990 640.240 1189.955 642.920 ;
        RECT 4.400 638.840 1189.955 640.240 ;
        RECT 3.990 630.720 1189.955 638.840 ;
        RECT 3.990 629.320 1189.070 630.720 ;
        RECT 3.990 626.640 1189.955 629.320 ;
        RECT 4.400 625.240 1189.955 626.640 ;
        RECT 3.990 617.120 1189.955 625.240 ;
        RECT 3.990 615.720 1189.070 617.120 ;
        RECT 3.990 613.040 1189.955 615.720 ;
        RECT 4.400 611.640 1189.955 613.040 ;
        RECT 3.990 604.880 1189.955 611.640 ;
        RECT 3.990 603.480 1189.070 604.880 ;
        RECT 3.990 599.440 1189.955 603.480 ;
        RECT 4.400 598.040 1189.955 599.440 ;
        RECT 3.990 591.280 1189.955 598.040 ;
        RECT 3.990 589.880 1189.070 591.280 ;
        RECT 3.990 587.200 1189.955 589.880 ;
        RECT 4.400 585.800 1189.955 587.200 ;
        RECT 3.990 577.680 1189.955 585.800 ;
        RECT 3.990 576.280 1189.070 577.680 ;
        RECT 3.990 573.600 1189.955 576.280 ;
        RECT 4.400 572.200 1189.955 573.600 ;
        RECT 3.990 564.080 1189.955 572.200 ;
        RECT 3.990 562.680 1189.070 564.080 ;
        RECT 3.990 560.000 1189.955 562.680 ;
        RECT 4.400 558.600 1189.955 560.000 ;
        RECT 3.990 550.480 1189.955 558.600 ;
        RECT 3.990 549.080 1189.070 550.480 ;
        RECT 3.990 546.400 1189.955 549.080 ;
        RECT 4.400 545.000 1189.955 546.400 ;
        RECT 3.990 536.880 1189.955 545.000 ;
        RECT 3.990 535.480 1189.070 536.880 ;
        RECT 3.990 532.800 1189.955 535.480 ;
        RECT 4.400 531.400 1189.955 532.800 ;
        RECT 3.990 523.280 1189.955 531.400 ;
        RECT 3.990 521.880 1189.070 523.280 ;
        RECT 3.990 519.200 1189.955 521.880 ;
        RECT 4.400 517.800 1189.955 519.200 ;
        RECT 3.990 509.680 1189.955 517.800 ;
        RECT 3.990 508.280 1189.070 509.680 ;
        RECT 3.990 505.600 1189.955 508.280 ;
        RECT 4.400 504.200 1189.955 505.600 ;
        RECT 3.990 496.080 1189.955 504.200 ;
        RECT 3.990 494.680 1189.070 496.080 ;
        RECT 3.990 492.000 1189.955 494.680 ;
        RECT 4.400 490.600 1189.955 492.000 ;
        RECT 3.990 482.480 1189.955 490.600 ;
        RECT 3.990 481.080 1189.070 482.480 ;
        RECT 3.990 478.400 1189.955 481.080 ;
        RECT 4.400 477.000 1189.955 478.400 ;
        RECT 3.990 468.880 1189.955 477.000 ;
        RECT 3.990 467.480 1189.070 468.880 ;
        RECT 3.990 464.800 1189.955 467.480 ;
        RECT 4.400 463.400 1189.955 464.800 ;
        RECT 3.990 455.280 1189.955 463.400 ;
        RECT 3.990 453.880 1189.070 455.280 ;
        RECT 3.990 451.200 1189.955 453.880 ;
        RECT 4.400 449.800 1189.955 451.200 ;
        RECT 3.990 441.680 1189.955 449.800 ;
        RECT 3.990 440.280 1189.070 441.680 ;
        RECT 3.990 437.600 1189.955 440.280 ;
        RECT 4.400 436.200 1189.955 437.600 ;
        RECT 3.990 428.080 1189.955 436.200 ;
        RECT 3.990 426.680 1189.070 428.080 ;
        RECT 3.990 424.000 1189.955 426.680 ;
        RECT 4.400 422.600 1189.955 424.000 ;
        RECT 3.990 414.480 1189.955 422.600 ;
        RECT 3.990 413.080 1189.070 414.480 ;
        RECT 3.990 410.400 1189.955 413.080 ;
        RECT 4.400 409.000 1189.955 410.400 ;
        RECT 3.990 400.880 1189.955 409.000 ;
        RECT 3.990 399.480 1189.070 400.880 ;
        RECT 3.990 396.800 1189.955 399.480 ;
        RECT 4.400 395.400 1189.955 396.800 ;
        RECT 3.990 387.280 1189.955 395.400 ;
        RECT 3.990 385.880 1189.070 387.280 ;
        RECT 3.990 383.200 1189.955 385.880 ;
        RECT 4.400 381.800 1189.955 383.200 ;
        RECT 3.990 373.680 1189.955 381.800 ;
        RECT 3.990 372.280 1189.070 373.680 ;
        RECT 3.990 369.600 1189.955 372.280 ;
        RECT 4.400 368.200 1189.955 369.600 ;
        RECT 3.990 360.080 1189.955 368.200 ;
        RECT 3.990 358.680 1189.070 360.080 ;
        RECT 3.990 356.000 1189.955 358.680 ;
        RECT 4.400 354.600 1189.955 356.000 ;
        RECT 3.990 346.480 1189.955 354.600 ;
        RECT 3.990 345.080 1189.070 346.480 ;
        RECT 3.990 342.400 1189.955 345.080 ;
        RECT 4.400 341.000 1189.955 342.400 ;
        RECT 3.990 332.880 1189.955 341.000 ;
        RECT 3.990 331.480 1189.070 332.880 ;
        RECT 3.990 328.800 1189.955 331.480 ;
        RECT 4.400 327.400 1189.955 328.800 ;
        RECT 3.990 319.280 1189.955 327.400 ;
        RECT 3.990 317.880 1189.070 319.280 ;
        RECT 3.990 315.200 1189.955 317.880 ;
        RECT 4.400 313.800 1189.955 315.200 ;
        RECT 3.990 307.040 1189.955 313.800 ;
        RECT 3.990 305.640 1189.070 307.040 ;
        RECT 3.990 301.600 1189.955 305.640 ;
        RECT 4.400 300.200 1189.955 301.600 ;
        RECT 3.990 293.440 1189.955 300.200 ;
        RECT 3.990 292.040 1189.070 293.440 ;
        RECT 3.990 289.360 1189.955 292.040 ;
        RECT 4.400 287.960 1189.955 289.360 ;
        RECT 3.990 279.840 1189.955 287.960 ;
        RECT 3.990 278.440 1189.070 279.840 ;
        RECT 3.990 275.760 1189.955 278.440 ;
        RECT 4.400 274.360 1189.955 275.760 ;
        RECT 3.990 266.240 1189.955 274.360 ;
        RECT 3.990 264.840 1189.070 266.240 ;
        RECT 3.990 262.160 1189.955 264.840 ;
        RECT 4.400 260.760 1189.955 262.160 ;
        RECT 3.990 252.640 1189.955 260.760 ;
        RECT 3.990 251.240 1189.070 252.640 ;
        RECT 3.990 248.560 1189.955 251.240 ;
        RECT 4.400 247.160 1189.955 248.560 ;
        RECT 3.990 239.040 1189.955 247.160 ;
        RECT 3.990 237.640 1189.070 239.040 ;
        RECT 3.990 234.960 1189.955 237.640 ;
        RECT 4.400 233.560 1189.955 234.960 ;
        RECT 3.990 225.440 1189.955 233.560 ;
        RECT 3.990 224.040 1189.070 225.440 ;
        RECT 3.990 221.360 1189.955 224.040 ;
        RECT 4.400 219.960 1189.955 221.360 ;
        RECT 3.990 211.840 1189.955 219.960 ;
        RECT 3.990 210.440 1189.070 211.840 ;
        RECT 3.990 207.760 1189.955 210.440 ;
        RECT 4.400 206.360 1189.955 207.760 ;
        RECT 3.990 198.240 1189.955 206.360 ;
        RECT 3.990 196.840 1189.070 198.240 ;
        RECT 3.990 194.160 1189.955 196.840 ;
        RECT 4.400 192.760 1189.955 194.160 ;
        RECT 3.990 184.640 1189.955 192.760 ;
        RECT 3.990 183.240 1189.070 184.640 ;
        RECT 3.990 180.560 1189.955 183.240 ;
        RECT 4.400 179.160 1189.955 180.560 ;
        RECT 3.990 171.040 1189.955 179.160 ;
        RECT 3.990 169.640 1189.070 171.040 ;
        RECT 3.990 166.960 1189.955 169.640 ;
        RECT 4.400 165.560 1189.955 166.960 ;
        RECT 3.990 157.440 1189.955 165.560 ;
        RECT 3.990 156.040 1189.070 157.440 ;
        RECT 3.990 153.360 1189.955 156.040 ;
        RECT 4.400 151.960 1189.955 153.360 ;
        RECT 3.990 143.840 1189.955 151.960 ;
        RECT 3.990 142.440 1189.070 143.840 ;
        RECT 3.990 139.760 1189.955 142.440 ;
        RECT 4.400 138.360 1189.955 139.760 ;
        RECT 3.990 130.240 1189.955 138.360 ;
        RECT 3.990 128.840 1189.070 130.240 ;
        RECT 3.990 126.160 1189.955 128.840 ;
        RECT 4.400 124.760 1189.955 126.160 ;
        RECT 3.990 116.640 1189.955 124.760 ;
        RECT 3.990 115.240 1189.070 116.640 ;
        RECT 3.990 112.560 1189.955 115.240 ;
        RECT 4.400 111.160 1189.955 112.560 ;
        RECT 3.990 103.040 1189.955 111.160 ;
        RECT 3.990 101.640 1189.070 103.040 ;
        RECT 3.990 98.960 1189.955 101.640 ;
        RECT 4.400 97.560 1189.955 98.960 ;
        RECT 3.990 89.440 1189.955 97.560 ;
        RECT 3.990 88.040 1189.070 89.440 ;
        RECT 3.990 85.360 1189.955 88.040 ;
        RECT 4.400 83.960 1189.955 85.360 ;
        RECT 3.990 75.840 1189.955 83.960 ;
        RECT 3.990 74.440 1189.070 75.840 ;
        RECT 3.990 71.760 1189.955 74.440 ;
        RECT 4.400 70.360 1189.955 71.760 ;
        RECT 3.990 62.240 1189.955 70.360 ;
        RECT 3.990 60.840 1189.070 62.240 ;
        RECT 3.990 58.160 1189.955 60.840 ;
        RECT 4.400 56.760 1189.955 58.160 ;
        RECT 3.990 48.640 1189.955 56.760 ;
        RECT 3.990 47.240 1189.070 48.640 ;
        RECT 3.990 44.560 1189.955 47.240 ;
        RECT 4.400 43.160 1189.955 44.560 ;
        RECT 3.990 35.040 1189.955 43.160 ;
        RECT 3.990 33.640 1189.070 35.040 ;
        RECT 3.990 30.960 1189.955 33.640 ;
        RECT 4.400 29.560 1189.955 30.960 ;
        RECT 3.990 21.440 1189.955 29.560 ;
        RECT 3.990 20.040 1189.070 21.440 ;
        RECT 3.990 17.360 1189.955 20.040 ;
        RECT 4.400 15.960 1189.955 17.360 ;
        RECT 3.990 9.200 1189.955 15.960 ;
        RECT 3.990 8.335 1189.070 9.200 ;
      LAYER met4 ;
        RECT 13.175 10.640 20.640 1191.600 ;
        RECT 23.040 10.640 97.440 1191.600 ;
        RECT 99.840 10.640 1174.640 1191.600 ;
  END
END register_file_16_1489f923c4dca729178b3e3233458550d8dddf29
END LIBRARY

