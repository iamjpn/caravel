magic
tech sky130A
magscale 1 2
timestamp 1607831768
<< obsli1 >>
rect 1104 2159 338836 177361
<< obsm1 >>
rect 1104 1776 338836 177472
<< metal2 >>
rect 5262 179200 5318 180000
rect 15842 179200 15898 180000
rect 26514 179200 26570 180000
rect 37094 179200 37150 180000
rect 47766 179200 47822 180000
rect 58346 179200 58402 180000
rect 69018 179200 69074 180000
rect 79598 179200 79654 180000
rect 90270 179200 90326 180000
rect 100850 179200 100906 180000
rect 111522 179200 111578 180000
rect 122102 179200 122158 180000
rect 132774 179200 132830 180000
rect 143354 179200 143410 180000
rect 154026 179200 154082 180000
rect 164606 179200 164662 180000
rect 175278 179200 175334 180000
rect 185858 179200 185914 180000
rect 196530 179200 196586 180000
rect 207110 179200 207166 180000
rect 217782 179200 217838 180000
rect 228362 179200 228418 180000
rect 239034 179200 239090 180000
rect 249614 179200 249670 180000
rect 260286 179200 260342 180000
rect 270866 179200 270922 180000
rect 281538 179200 281594 180000
rect 292118 179200 292174 180000
rect 302790 179200 302846 180000
rect 313370 179200 313426 180000
rect 324042 179200 324098 180000
rect 334622 179200 334678 180000
rect 5262 0 5318 800
rect 15842 0 15898 800
rect 26514 0 26570 800
rect 37094 0 37150 800
rect 47766 0 47822 800
rect 58346 0 58402 800
rect 69018 0 69074 800
rect 79598 0 79654 800
rect 90270 0 90326 800
rect 100850 0 100906 800
rect 111522 0 111578 800
rect 122102 0 122158 800
rect 132774 0 132830 800
rect 143354 0 143410 800
rect 154026 0 154082 800
rect 164606 0 164662 800
rect 175278 0 175334 800
rect 185858 0 185914 800
rect 196530 0 196586 800
rect 207110 0 207166 800
rect 217782 0 217838 800
rect 228362 0 228418 800
rect 239034 0 239090 800
rect 249614 0 249670 800
rect 260286 0 260342 800
rect 270866 0 270922 800
rect 281538 0 281594 800
rect 292118 0 292174 800
rect 302790 0 302846 800
rect 313370 0 313426 800
rect 324042 0 324098 800
rect 334622 0 334678 800
<< obsm2 >>
rect 1400 179144 5206 179200
rect 5374 179144 15786 179200
rect 15954 179144 26458 179200
rect 26626 179144 37038 179200
rect 37206 179144 47710 179200
rect 47878 179144 58290 179200
rect 58458 179144 68962 179200
rect 69130 179144 79542 179200
rect 79710 179144 90214 179200
rect 90382 179144 100794 179200
rect 100962 179144 111466 179200
rect 111634 179144 122046 179200
rect 122214 179144 132718 179200
rect 132886 179144 143298 179200
rect 143466 179144 153970 179200
rect 154138 179144 164550 179200
rect 164718 179144 175222 179200
rect 175390 179144 185802 179200
rect 185970 179144 196474 179200
rect 196642 179144 207054 179200
rect 207222 179144 217726 179200
rect 217894 179144 228306 179200
rect 228474 179144 238978 179200
rect 239146 179144 249558 179200
rect 249726 179144 260230 179200
rect 260398 179144 270810 179200
rect 270978 179144 281482 179200
rect 281650 179144 292062 179200
rect 292230 179144 302734 179200
rect 302902 179144 313314 179200
rect 313482 179144 323986 179200
rect 324154 179144 334566 179200
rect 334734 179144 338264 179200
rect 1400 856 338264 179144
rect 1400 800 5206 856
rect 5374 800 15786 856
rect 15954 800 26458 856
rect 26626 800 37038 856
rect 37206 800 47710 856
rect 47878 800 58290 856
rect 58458 800 68962 856
rect 69130 800 79542 856
rect 79710 800 90214 856
rect 90382 800 100794 856
rect 100962 800 111466 856
rect 111634 800 122046 856
rect 122214 800 132718 856
rect 132886 800 143298 856
rect 143466 800 153970 856
rect 154138 800 164550 856
rect 164718 800 175222 856
rect 175390 800 185802 856
rect 185970 800 196474 856
rect 196642 800 207054 856
rect 207222 800 217726 856
rect 217894 800 228306 856
rect 228474 800 238978 856
rect 239146 800 249558 856
rect 249726 800 260230 856
rect 260398 800 270810 856
rect 270978 800 281482 856
rect 281650 800 292062 856
rect 292230 800 302734 856
rect 302902 800 313314 856
rect 313482 800 323986 856
rect 324154 800 334566 856
rect 334734 800 338264 856
<< metal3 >>
rect 0 174360 800 174480
rect 0 163072 800 163192
rect 0 151784 800 151904
rect 0 140632 800 140752
rect 0 129344 800 129464
rect 0 118056 800 118176
rect 0 106768 800 106888
rect 0 95616 800 95736
rect 0 84328 800 84448
rect 0 73040 800 73160
rect 0 61752 800 61872
rect 0 50600 800 50720
rect 0 39312 800 39432
rect 0 28024 800 28144
rect 0 16736 800 16856
rect 0 5584 800 5704
<< obsm3 >>
rect 800 174560 337259 177377
rect 880 174280 337259 174560
rect 800 163272 337259 174280
rect 880 162992 337259 163272
rect 800 151984 337259 162992
rect 880 151704 337259 151984
rect 800 140832 337259 151704
rect 880 140552 337259 140832
rect 800 129544 337259 140552
rect 880 129264 337259 129544
rect 800 118256 337259 129264
rect 880 117976 337259 118256
rect 800 106968 337259 117976
rect 880 106688 337259 106968
rect 800 95816 337259 106688
rect 880 95536 337259 95816
rect 800 84528 337259 95536
rect 880 84248 337259 84528
rect 800 73240 337259 84248
rect 880 72960 337259 73240
rect 800 61952 337259 72960
rect 880 61672 337259 61952
rect 800 50800 337259 61672
rect 880 50520 337259 50800
rect 800 39512 337259 50520
rect 880 39232 337259 39512
rect 800 28224 337259 39232
rect 880 27944 337259 28224
rect 800 16936 337259 27944
rect 880 16656 337259 16936
rect 800 5784 337259 16656
rect 880 5504 337259 5784
rect 800 2143 337259 5504
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
<< obsm4 >>
rect 5947 2128 19488 177392
rect 19968 2128 335005 177392
<< obsm5 >>
rect 230300 47100 281404 101140
<< labels >>
rlabel metal3 s 0 5584 800 5704 6 A[0]
port 1 nsew default input
rlabel metal3 s 0 16736 800 16856 6 A[1]
port 2 nsew default input
rlabel metal3 s 0 28024 800 28144 6 A[2]
port 3 nsew default input
rlabel metal3 s 0 39312 800 39432 6 A[3]
port 4 nsew default input
rlabel metal3 s 0 50600 800 50720 6 A[4]
port 5 nsew default input
rlabel metal3 s 0 61752 800 61872 6 A[5]
port 6 nsew default input
rlabel metal3 s 0 73040 800 73160 6 A[6]
port 7 nsew default input
rlabel metal3 s 0 84328 800 84448 6 A[7]
port 8 nsew default input
rlabel metal3 s 0 95616 800 95736 6 A[8]
port 9 nsew default input
rlabel metal3 s 0 106768 800 106888 6 A[9]
port 10 nsew default input
rlabel metal3 s 0 118056 800 118176 6 CLK
port 11 nsew default input
rlabel metal2 s 5262 179200 5318 180000 6 Di[0]
port 12 nsew default input
rlabel metal2 s 111522 179200 111578 180000 6 Di[10]
port 13 nsew default input
rlabel metal2 s 122102 179200 122158 180000 6 Di[11]
port 14 nsew default input
rlabel metal2 s 132774 179200 132830 180000 6 Di[12]
port 15 nsew default input
rlabel metal2 s 143354 179200 143410 180000 6 Di[13]
port 16 nsew default input
rlabel metal2 s 154026 179200 154082 180000 6 Di[14]
port 17 nsew default input
rlabel metal2 s 164606 179200 164662 180000 6 Di[15]
port 18 nsew default input
rlabel metal2 s 175278 179200 175334 180000 6 Di[16]
port 19 nsew default input
rlabel metal2 s 185858 179200 185914 180000 6 Di[17]
port 20 nsew default input
rlabel metal2 s 196530 179200 196586 180000 6 Di[18]
port 21 nsew default input
rlabel metal2 s 207110 179200 207166 180000 6 Di[19]
port 22 nsew default input
rlabel metal2 s 15842 179200 15898 180000 6 Di[1]
port 23 nsew default input
rlabel metal2 s 217782 179200 217838 180000 6 Di[20]
port 24 nsew default input
rlabel metal2 s 228362 179200 228418 180000 6 Di[21]
port 25 nsew default input
rlabel metal2 s 239034 179200 239090 180000 6 Di[22]
port 26 nsew default input
rlabel metal2 s 249614 179200 249670 180000 6 Di[23]
port 27 nsew default input
rlabel metal2 s 260286 179200 260342 180000 6 Di[24]
port 28 nsew default input
rlabel metal2 s 270866 179200 270922 180000 6 Di[25]
port 29 nsew default input
rlabel metal2 s 281538 179200 281594 180000 6 Di[26]
port 30 nsew default input
rlabel metal2 s 292118 179200 292174 180000 6 Di[27]
port 31 nsew default input
rlabel metal2 s 302790 179200 302846 180000 6 Di[28]
port 32 nsew default input
rlabel metal2 s 313370 179200 313426 180000 6 Di[29]
port 33 nsew default input
rlabel metal2 s 26514 179200 26570 180000 6 Di[2]
port 34 nsew default input
rlabel metal2 s 324042 179200 324098 180000 6 Di[30]
port 35 nsew default input
rlabel metal2 s 334622 179200 334678 180000 6 Di[31]
port 36 nsew default input
rlabel metal2 s 37094 179200 37150 180000 6 Di[3]
port 37 nsew default input
rlabel metal2 s 47766 179200 47822 180000 6 Di[4]
port 38 nsew default input
rlabel metal2 s 58346 179200 58402 180000 6 Di[5]
port 39 nsew default input
rlabel metal2 s 69018 179200 69074 180000 6 Di[6]
port 40 nsew default input
rlabel metal2 s 79598 179200 79654 180000 6 Di[7]
port 41 nsew default input
rlabel metal2 s 90270 179200 90326 180000 6 Di[8]
port 42 nsew default input
rlabel metal2 s 100850 179200 100906 180000 6 Di[9]
port 43 nsew default input
rlabel metal2 s 5262 0 5318 800 6 Do[0]
port 44 nsew default output
rlabel metal2 s 111522 0 111578 800 6 Do[10]
port 45 nsew default output
rlabel metal2 s 122102 0 122158 800 6 Do[11]
port 46 nsew default output
rlabel metal2 s 132774 0 132830 800 6 Do[12]
port 47 nsew default output
rlabel metal2 s 143354 0 143410 800 6 Do[13]
port 48 nsew default output
rlabel metal2 s 154026 0 154082 800 6 Do[14]
port 49 nsew default output
rlabel metal2 s 164606 0 164662 800 6 Do[15]
port 50 nsew default output
rlabel metal2 s 175278 0 175334 800 6 Do[16]
port 51 nsew default output
rlabel metal2 s 185858 0 185914 800 6 Do[17]
port 52 nsew default output
rlabel metal2 s 196530 0 196586 800 6 Do[18]
port 53 nsew default output
rlabel metal2 s 207110 0 207166 800 6 Do[19]
port 54 nsew default output
rlabel metal2 s 15842 0 15898 800 6 Do[1]
port 55 nsew default output
rlabel metal2 s 217782 0 217838 800 6 Do[20]
port 56 nsew default output
rlabel metal2 s 228362 0 228418 800 6 Do[21]
port 57 nsew default output
rlabel metal2 s 239034 0 239090 800 6 Do[22]
port 58 nsew default output
rlabel metal2 s 249614 0 249670 800 6 Do[23]
port 59 nsew default output
rlabel metal2 s 260286 0 260342 800 6 Do[24]
port 60 nsew default output
rlabel metal2 s 270866 0 270922 800 6 Do[25]
port 61 nsew default output
rlabel metal2 s 281538 0 281594 800 6 Do[26]
port 62 nsew default output
rlabel metal2 s 292118 0 292174 800 6 Do[27]
port 63 nsew default output
rlabel metal2 s 302790 0 302846 800 6 Do[28]
port 64 nsew default output
rlabel metal2 s 313370 0 313426 800 6 Do[29]
port 65 nsew default output
rlabel metal2 s 26514 0 26570 800 6 Do[2]
port 66 nsew default output
rlabel metal2 s 324042 0 324098 800 6 Do[30]
port 67 nsew default output
rlabel metal2 s 334622 0 334678 800 6 Do[31]
port 68 nsew default output
rlabel metal2 s 37094 0 37150 800 6 Do[3]
port 69 nsew default output
rlabel metal2 s 47766 0 47822 800 6 Do[4]
port 70 nsew default output
rlabel metal2 s 58346 0 58402 800 6 Do[5]
port 71 nsew default output
rlabel metal2 s 69018 0 69074 800 6 Do[6]
port 72 nsew default output
rlabel metal2 s 79598 0 79654 800 6 Do[7]
port 73 nsew default output
rlabel metal2 s 90270 0 90326 800 6 Do[8]
port 74 nsew default output
rlabel metal2 s 100850 0 100906 800 6 Do[9]
port 75 nsew default output
rlabel metal3 s 0 174360 800 174480 6 EN
port 76 nsew default input
rlabel metal3 s 0 129344 800 129464 6 WE[0]
port 77 nsew default input
rlabel metal3 s 0 140632 800 140752 6 WE[1]
port 78 nsew default input
rlabel metal3 s 0 151784 800 151904 6 WE[2]
port 79 nsew default input
rlabel metal3 s 0 163072 800 163192 6 WE[3]
port 80 nsew default input
rlabel metal4 s 4208 2128 4528 177392 6 VPWR
port 81 nsew power input
rlabel metal4 s 19568 2128 19888 177392 6 VGND
port 82 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 338874 180000
string LEFview TRUE
<< end >>
