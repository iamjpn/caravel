module register_file_16_1489f923c4dca729178b3e3233458550d8dddf29(clk, d_in, w_in, dbg_gpr_req, dbg_gpr_addr, sim_dump, d_out, dbg_gpr_ack, dbg_gpr_data, sim_dump_done, log_out);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire [6:0] _04_;
  wire _05_;
  wire [63:0] _06_;
  wire _07_;
  wire [63:0] _08_;
  wire _09_;
  wire [63:0] _10_;
  wire [191:0] _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire [63:0] _18_;
  wire [8191:0] _19_;
  wire [63:0] _20_;
  wire [8191:0] _21_;
  wire [8191:0] _22_;
  wire [63:0] _23_;
  input clk;
  input [23:0] d_in;
  output [191:0] d_out;
  reg dbg_ack;
  reg [63:0] dbg_data;
  output dbg_gpr_ack;
  input [6:0] dbg_gpr_addr;
  output [63:0] dbg_gpr_data;
  input dbg_gpr_req;
  output [71:0] log_out;
  wire [63:0] rd_port_b;
  reg [71:0] \rf_log.log_data ;
  input sim_dump;
  output sim_dump_done;
  input [71:0] w_in;
  reg [63:0] \$mem$\10022  [127:0];
  reg [63:0] \10022  [127:0];
  initial begin
    \10022 [0] = 64'h0000000000000000;
    \10022 [1] = 64'h0000000000000000;
    \10022 [2] = 64'h0000000000000000;
    \10022 [3] = 64'h0000000000000000;
    \10022 [4] = 64'h0000000000000000;
    \10022 [5] = 64'h0000000000000000;
    \10022 [6] = 64'h0000000000000000;
    \10022 [7] = 64'h0000000000000000;
    \10022 [8] = 64'h0000000000000000;
    \10022 [9] = 64'h0000000000000000;
    \10022 [10] = 64'h0000000000000000;
    \10022 [11] = 64'h0000000000000000;
    \10022 [12] = 64'h0000000000000000;
    \10022 [13] = 64'h0000000000000000;
    \10022 [14] = 64'h0000000000000000;
    \10022 [15] = 64'h0000000000000000;
    \10022 [16] = 64'h0000000000000000;
    \10022 [17] = 64'h0000000000000000;
    \10022 [18] = 64'h0000000000000000;
    \10022 [19] = 64'h0000000000000000;
    \10022 [20] = 64'h0000000000000000;
    \10022 [21] = 64'h0000000000000000;
    \10022 [22] = 64'h0000000000000000;
    \10022 [23] = 64'h0000000000000000;
    \10022 [24] = 64'h0000000000000000;
    \10022 [25] = 64'h0000000000000000;
    \10022 [26] = 64'h0000000000000000;
    \10022 [27] = 64'h0000000000000000;
    \10022 [28] = 64'h0000000000000000;
    \10022 [29] = 64'h0000000000000000;
    \10022 [30] = 64'h0000000000000000;
    \10022 [31] = 64'h0000000000000000;
    \10022 [32] = 64'h0000000000000000;
    \10022 [33] = 64'h0000000000000000;
    \10022 [34] = 64'h0000000000000000;
    \10022 [35] = 64'h0000000000000000;
    \10022 [36] = 64'h0000000000000000;
    \10022 [37] = 64'h0000000000000000;
    \10022 [38] = 64'h0000000000000000;
    \10022 [39] = 64'h0000000000000000;
    \10022 [40] = 64'h0000000000000000;
    \10022 [41] = 64'h0000000000000000;
    \10022 [42] = 64'h0000000000000000;
    \10022 [43] = 64'h0000000000000000;
    \10022 [44] = 64'h0000000000000000;
    \10022 [45] = 64'h0000000000000000;
    \10022 [46] = 64'h0000000000000000;
    \10022 [47] = 64'h0000000000000000;
    \10022 [48] = 64'h0000000000000000;
    \10022 [49] = 64'h0000000000000000;
    \10022 [50] = 64'h0000000000000000;
    \10022 [51] = 64'h0000000000000000;
    \10022 [52] = 64'h0000000000000000;
    \10022 [53] = 64'h0000000000000000;
    \10022 [54] = 64'h0000000000000000;
    \10022 [55] = 64'h0000000000000000;
    \10022 [56] = 64'h0000000000000000;
    \10022 [57] = 64'h0000000000000000;
    \10022 [58] = 64'h0000000000000000;
    \10022 [59] = 64'h0000000000000000;
    \10022 [60] = 64'h0000000000000000;
    \10022 [61] = 64'h0000000000000000;
    \10022 [62] = 64'h0000000000000000;
    \10022 [63] = 64'h0000000000000000;
    \10022 [64] = 64'h0000000000000000;
    \10022 [65] = 64'h0000000000000000;
    \10022 [66] = 64'h0000000000000000;
    \10022 [67] = 64'h0000000000000000;
    \10022 [68] = 64'h0000000000000000;
    \10022 [69] = 64'h0000000000000000;
    \10022 [70] = 64'h0000000000000000;
    \10022 [71] = 64'h0000000000000000;
    \10022 [72] = 64'h0000000000000000;
    \10022 [73] = 64'h0000000000000000;
    \10022 [74] = 64'h0000000000000000;
    \10022 [75] = 64'h0000000000000000;
    \10022 [76] = 64'h0000000000000000;
    \10022 [77] = 64'h0000000000000000;
    \10022 [78] = 64'h0000000000000000;
    \10022 [79] = 64'h0000000000000000;
    \10022 [80] = 64'h0000000000000000;
    \10022 [81] = 64'h0000000000000000;
    \10022 [82] = 64'h0000000000000000;
    \10022 [83] = 64'h0000000000000000;
    \10022 [84] = 64'h0000000000000000;
    \10022 [85] = 64'h0000000000000000;
    \10022 [86] = 64'h0000000000000000;
    \10022 [87] = 64'h0000000000000000;
    \10022 [88] = 64'h0000000000000000;
    \10022 [89] = 64'h0000000000000000;
    \10022 [90] = 64'h0000000000000000;
    \10022 [91] = 64'h0000000000000000;
    \10022 [92] = 64'h0000000000000000;
    \10022 [93] = 64'h0000000000000000;
    \10022 [94] = 64'h0000000000000000;
    \10022 [95] = 64'h0000000000000000;
    \10022 [96] = 64'h0000000000000000;
    \10022 [97] = 64'h0000000000000000;
    \10022 [98] = 64'h0000000000000000;
    \10022 [99] = 64'h0000000000000000;
    \10022 [100] = 64'h0000000000000000;
    \10022 [101] = 64'h0000000000000000;
    \10022 [102] = 64'h0000000000000000;
    \10022 [103] = 64'h0000000000000000;
    \10022 [104] = 64'h0000000000000000;
    \10022 [105] = 64'h0000000000000000;
    \10022 [106] = 64'h0000000000000000;
    \10022 [107] = 64'h0000000000000000;
    \10022 [108] = 64'h0000000000000000;
    \10022 [109] = 64'h0000000000000000;
    \10022 [110] = 64'h0000000000000000;
    \10022 [111] = 64'h0000000000000000;
    \10022 [112] = 64'h0000000000000000;
    \10022 [113] = 64'h0000000000000000;
    \10022 [114] = 64'h0000000000000000;
    \10022 [115] = 64'h0000000000000000;
    \10022 [116] = 64'h0000000000000000;
    \10022 [117] = 64'h0000000000000000;
    \10022 [118] = 64'h0000000000000000;
    \10022 [119] = 64'h0000000000000000;
    \10022 [120] = 64'h0000000000000000;
    \10022 [121] = 64'h0000000000000000;
    \10022 [122] = 64'h0000000000000000;
    \10022 [123] = 64'h0000000000000000;
    \10022 [124] = 64'h0000000000000000;
    \10022 [125] = 64'h0000000000000000;
    \10022 [126] = 64'h0000000000000000;
    \10022 [127] = 64'h0000000000000000;
  end
  always @(posedge clk) begin
    if (w_in[71]) \10022 [{ 1'h0, w_in[5:0] }] <= w_in[70:7];
  end
  assign _20_ = \10022 [{ 1'h0, d_in[22:17] }];
  assign rd_port_b = \10022 [_04_];
  assign _23_ = \10022 [{ 1'h0, d_in[6:1] }];
  assign _17_ = dbg_gpr_req ? _15_ : 1'h0;
  assign _18_ = _16_ ? rd_port_b : dbg_data;
  always @(posedge clk)
    dbg_data <= _18_;
  always @(posedge clk)
    dbg_ack <= _17_;
  always @(posedge clk)
    \rf_log.log_data  <= { w_in[70:7], w_in[71], w_in[6:0] };
  assign _00_ = ~ d_in[8];
  assign _01_ = _00_ & dbg_gpr_req;
  assign _02_ = ~ dbg_ack;
  assign _03_ = _01_ & _02_;
  assign _04_ = _03_ ? { 1'h0, dbg_gpr_addr[5:0] } : { 1'h0, d_in[14:9] };
  assign _05_ = { 1'h0, d_in[6:1] } == { 1'h0, w_in[5:0] };
  assign _06_ = _05_ ? w_in[70:7] : _23_;
  assign _07_ = _04_ == { 1'h0, w_in[5:0] };
  assign _08_ = _07_ ? w_in[70:7] : rd_port_b;
  assign _09_ = { 1'h0, d_in[22:17] } == { 1'h0, w_in[5:0] };
  assign _10_ = _09_ ? w_in[70:7] : _20_;
  assign _11_ = w_in[71] ? { _10_, _08_, _06_ } : { _20_, rd_port_b, _23_ };
  assign _12_ = ~ d_in[8];
  assign _13_ = ~ dbg_ack;
  assign _14_ = _12_ & _13_;
  assign _15_ = _14_ ? 1'h1 : dbg_ack;
  assign _16_ = dbg_gpr_req & _14_;
  assign d_out = _11_;
  assign dbg_gpr_ack = dbg_ack;
  assign dbg_gpr_data = dbg_data;
  assign sim_dump_done = 1'h0;
  assign log_out = \rf_log.log_data ;
endmodule
