magic
tech sky130A
magscale 1 2
timestamp 1607842331
<< obsli1 >>
rect 1104 2159 237544 238289
<< obsm1 >>
rect 566 892 237544 238740
<< metal2 >>
rect 1674 240038 1730 240838
rect 3514 240038 3570 240838
rect 5354 240038 5410 240838
rect 7194 240038 7250 240838
rect 9034 240038 9090 240838
rect 10874 240038 10930 240838
rect 12714 240038 12770 240838
rect 14554 240038 14610 240838
rect 16394 240038 16450 240838
rect 18234 240038 18290 240838
rect 20074 240038 20130 240838
rect 21914 240038 21970 240838
rect 23754 240038 23810 240838
rect 25594 240038 25650 240838
rect 27434 240038 27490 240838
rect 29274 240038 29330 240838
rect 31114 240038 31170 240838
rect 32954 240038 33010 240838
rect 34794 240038 34850 240838
rect 36634 240038 36690 240838
rect 38290 240038 38346 240838
rect 40130 240038 40186 240838
rect 41970 240038 42026 240838
rect 43810 240038 43866 240838
rect 45650 240038 45706 240838
rect 47490 240038 47546 240838
rect 49330 240038 49386 240838
rect 51170 240038 51226 240838
rect 53010 240038 53066 240838
rect 54850 240038 54906 240838
rect 56690 240038 56746 240838
rect 58530 240038 58586 240838
rect 60370 240038 60426 240838
rect 62210 240038 62266 240838
rect 64050 240038 64106 240838
rect 65890 240038 65946 240838
rect 67730 240038 67786 240838
rect 69570 240038 69626 240838
rect 71410 240038 71466 240838
rect 73250 240038 73306 240838
rect 75090 240038 75146 240838
rect 76930 240038 76986 240838
rect 78586 240038 78642 240838
rect 80426 240038 80482 240838
rect 82266 240038 82322 240838
rect 84106 240038 84162 240838
rect 85946 240038 86002 240838
rect 87786 240038 87842 240838
rect 89626 240038 89682 240838
rect 91466 240038 91522 240838
rect 93306 240038 93362 240838
rect 95146 240038 95202 240838
rect 96986 240038 97042 240838
rect 98826 240038 98882 240838
rect 100666 240038 100722 240838
rect 102506 240038 102562 240838
rect 104346 240038 104402 240838
rect 106186 240038 106242 240838
rect 108026 240038 108082 240838
rect 109866 240038 109922 240838
rect 111706 240038 111762 240838
rect 113546 240038 113602 240838
rect 115386 240038 115442 240838
rect 117226 240038 117282 240838
rect 118882 240038 118938 240838
rect 120722 240038 120778 240838
rect 122562 240038 122618 240838
rect 124402 240038 124458 240838
rect 126242 240038 126298 240838
rect 128082 240038 128138 240838
rect 129922 240038 129978 240838
rect 131762 240038 131818 240838
rect 133602 240038 133658 240838
rect 135442 240038 135498 240838
rect 137282 240038 137338 240838
rect 139122 240038 139178 240838
rect 140962 240038 141018 240838
rect 142802 240038 142858 240838
rect 144642 240038 144698 240838
rect 146482 240038 146538 240838
rect 148322 240038 148378 240838
rect 150162 240038 150218 240838
rect 152002 240038 152058 240838
rect 153842 240038 153898 240838
rect 155682 240038 155738 240838
rect 157522 240038 157578 240838
rect 159178 240038 159234 240838
rect 161018 240038 161074 240838
rect 162858 240038 162914 240838
rect 164698 240038 164754 240838
rect 166538 240038 166594 240838
rect 168378 240038 168434 240838
rect 170218 240038 170274 240838
rect 172058 240038 172114 240838
rect 173898 240038 173954 240838
rect 175738 240038 175794 240838
rect 177578 240038 177634 240838
rect 179418 240038 179474 240838
rect 181258 240038 181314 240838
rect 183098 240038 183154 240838
rect 184938 240038 184994 240838
rect 186778 240038 186834 240838
rect 188618 240038 188674 240838
rect 190458 240038 190514 240838
rect 192298 240038 192354 240838
rect 194138 240038 194194 240838
rect 195978 240038 196034 240838
rect 197818 240038 197874 240838
rect 199474 240038 199530 240838
rect 201314 240038 201370 240838
rect 203154 240038 203210 240838
rect 204994 240038 205050 240838
rect 206834 240038 206890 240838
rect 208674 240038 208730 240838
rect 210514 240038 210570 240838
rect 212354 240038 212410 240838
rect 214194 240038 214250 240838
rect 216034 240038 216090 240838
rect 217874 240038 217930 240838
rect 219714 240038 219770 240838
rect 221554 240038 221610 240838
rect 223394 240038 223450 240838
rect 225234 240038 225290 240838
rect 227074 240038 227130 240838
rect 228914 240038 228970 240838
rect 230754 240038 230810 240838
rect 232594 240038 232650 240838
rect 234434 240038 234490 240838
rect 236274 240038 236330 240838
rect 237930 240038 237986 240838
rect 570 0 626 800
rect 2226 0 2282 800
rect 4066 0 4122 800
rect 5906 0 5962 800
rect 7746 0 7802 800
rect 9586 0 9642 800
rect 11426 0 11482 800
rect 13266 0 13322 800
rect 15106 0 15162 800
rect 16946 0 17002 800
rect 18786 0 18842 800
rect 20626 0 20682 800
rect 22466 0 22522 800
rect 24306 0 24362 800
rect 26146 0 26202 800
rect 27986 0 28042 800
rect 29826 0 29882 800
rect 31666 0 31722 800
rect 33506 0 33562 800
rect 35346 0 35402 800
rect 37186 0 37242 800
rect 39026 0 39082 800
rect 40682 0 40738 800
rect 42522 0 42578 800
rect 44362 0 44418 800
rect 46202 0 46258 800
rect 48042 0 48098 800
rect 49882 0 49938 800
rect 51722 0 51778 800
rect 53562 0 53618 800
rect 55402 0 55458 800
rect 57242 0 57298 800
rect 59082 0 59138 800
rect 60922 0 60978 800
rect 62762 0 62818 800
rect 64602 0 64658 800
rect 66442 0 66498 800
rect 68282 0 68338 800
rect 70122 0 70178 800
rect 71962 0 72018 800
rect 73802 0 73858 800
rect 75642 0 75698 800
rect 77482 0 77538 800
rect 79322 0 79378 800
rect 80978 0 81034 800
rect 82818 0 82874 800
rect 84658 0 84714 800
rect 86498 0 86554 800
rect 88338 0 88394 800
rect 90178 0 90234 800
rect 92018 0 92074 800
rect 93858 0 93914 800
rect 95698 0 95754 800
rect 97538 0 97594 800
rect 99378 0 99434 800
rect 101218 0 101274 800
rect 103058 0 103114 800
rect 104898 0 104954 800
rect 106738 0 106794 800
rect 108578 0 108634 800
rect 110418 0 110474 800
rect 112258 0 112314 800
rect 114098 0 114154 800
rect 115938 0 115994 800
rect 117778 0 117834 800
rect 119618 0 119674 800
rect 121274 0 121330 800
rect 123114 0 123170 800
rect 124954 0 125010 800
rect 126794 0 126850 800
rect 128634 0 128690 800
rect 130474 0 130530 800
rect 132314 0 132370 800
rect 134154 0 134210 800
rect 135994 0 136050 800
rect 137834 0 137890 800
rect 139674 0 139730 800
rect 141514 0 141570 800
rect 143354 0 143410 800
rect 145194 0 145250 800
rect 147034 0 147090 800
rect 148874 0 148930 800
rect 150714 0 150770 800
rect 152554 0 152610 800
rect 154394 0 154450 800
rect 156234 0 156290 800
rect 158074 0 158130 800
rect 159914 0 159970 800
rect 161570 0 161626 800
rect 163410 0 163466 800
rect 165250 0 165306 800
rect 167090 0 167146 800
rect 168930 0 168986 800
rect 170770 0 170826 800
rect 172610 0 172666 800
rect 174450 0 174506 800
rect 176290 0 176346 800
rect 178130 0 178186 800
rect 179970 0 180026 800
rect 181810 0 181866 800
rect 183650 0 183706 800
rect 185490 0 185546 800
rect 187330 0 187386 800
rect 189170 0 189226 800
rect 191010 0 191066 800
rect 192850 0 192906 800
rect 194690 0 194746 800
rect 196530 0 196586 800
rect 198370 0 198426 800
rect 200210 0 200266 800
rect 201866 0 201922 800
rect 203706 0 203762 800
rect 205546 0 205602 800
rect 207386 0 207442 800
rect 209226 0 209282 800
rect 211066 0 211122 800
rect 212906 0 212962 800
rect 214746 0 214802 800
rect 216586 0 216642 800
rect 218426 0 218482 800
rect 220266 0 220322 800
rect 222106 0 222162 800
rect 223946 0 224002 800
rect 225786 0 225842 800
rect 227626 0 227682 800
rect 229466 0 229522 800
rect 231306 0 231362 800
rect 233146 0 233202 800
rect 234986 0 235042 800
rect 236826 0 236882 800
<< obsm2 >>
rect 572 239982 1618 240038
rect 1786 239982 3458 240038
rect 3626 239982 5298 240038
rect 5466 239982 7138 240038
rect 7306 239982 8978 240038
rect 9146 239982 10818 240038
rect 10986 239982 12658 240038
rect 12826 239982 14498 240038
rect 14666 239982 16338 240038
rect 16506 239982 18178 240038
rect 18346 239982 20018 240038
rect 20186 239982 21858 240038
rect 22026 239982 23698 240038
rect 23866 239982 25538 240038
rect 25706 239982 27378 240038
rect 27546 239982 29218 240038
rect 29386 239982 31058 240038
rect 31226 239982 32898 240038
rect 33066 239982 34738 240038
rect 34906 239982 36578 240038
rect 36746 239982 38234 240038
rect 38402 239982 40074 240038
rect 40242 239982 41914 240038
rect 42082 239982 43754 240038
rect 43922 239982 45594 240038
rect 45762 239982 47434 240038
rect 47602 239982 49274 240038
rect 49442 239982 51114 240038
rect 51282 239982 52954 240038
rect 53122 239982 54794 240038
rect 54962 239982 56634 240038
rect 56802 239982 58474 240038
rect 58642 239982 60314 240038
rect 60482 239982 62154 240038
rect 62322 239982 63994 240038
rect 64162 239982 65834 240038
rect 66002 239982 67674 240038
rect 67842 239982 69514 240038
rect 69682 239982 71354 240038
rect 71522 239982 73194 240038
rect 73362 239982 75034 240038
rect 75202 239982 76874 240038
rect 77042 239982 78530 240038
rect 78698 239982 80370 240038
rect 80538 239982 82210 240038
rect 82378 239982 84050 240038
rect 84218 239982 85890 240038
rect 86058 239982 87730 240038
rect 87898 239982 89570 240038
rect 89738 239982 91410 240038
rect 91578 239982 93250 240038
rect 93418 239982 95090 240038
rect 95258 239982 96930 240038
rect 97098 239982 98770 240038
rect 98938 239982 100610 240038
rect 100778 239982 102450 240038
rect 102618 239982 104290 240038
rect 104458 239982 106130 240038
rect 106298 239982 107970 240038
rect 108138 239982 109810 240038
rect 109978 239982 111650 240038
rect 111818 239982 113490 240038
rect 113658 239982 115330 240038
rect 115498 239982 117170 240038
rect 117338 239982 118826 240038
rect 118994 239982 120666 240038
rect 120834 239982 122506 240038
rect 122674 239982 124346 240038
rect 124514 239982 126186 240038
rect 126354 239982 128026 240038
rect 128194 239982 129866 240038
rect 130034 239982 131706 240038
rect 131874 239982 133546 240038
rect 133714 239982 135386 240038
rect 135554 239982 137226 240038
rect 137394 239982 139066 240038
rect 139234 239982 140906 240038
rect 141074 239982 142746 240038
rect 142914 239982 144586 240038
rect 144754 239982 146426 240038
rect 146594 239982 148266 240038
rect 148434 239982 150106 240038
rect 150274 239982 151946 240038
rect 152114 239982 153786 240038
rect 153954 239982 155626 240038
rect 155794 239982 157466 240038
rect 157634 239982 159122 240038
rect 159290 239982 160962 240038
rect 161130 239982 162802 240038
rect 162970 239982 164642 240038
rect 164810 239982 166482 240038
rect 166650 239982 168322 240038
rect 168490 239982 170162 240038
rect 170330 239982 172002 240038
rect 172170 239982 173842 240038
rect 174010 239982 175682 240038
rect 175850 239982 177522 240038
rect 177690 239982 179362 240038
rect 179530 239982 181202 240038
rect 181370 239982 183042 240038
rect 183210 239982 184882 240038
rect 185050 239982 186722 240038
rect 186890 239982 188562 240038
rect 188730 239982 190402 240038
rect 190570 239982 192242 240038
rect 192410 239982 194082 240038
rect 194250 239982 195922 240038
rect 196090 239982 197762 240038
rect 197930 239982 199418 240038
rect 199586 239982 201258 240038
rect 201426 239982 203098 240038
rect 203266 239982 204938 240038
rect 205106 239982 206778 240038
rect 206946 239982 208618 240038
rect 208786 239982 210458 240038
rect 210626 239982 212298 240038
rect 212466 239982 214138 240038
rect 214306 239982 215978 240038
rect 216146 239982 217818 240038
rect 217986 239982 219658 240038
rect 219826 239982 221498 240038
rect 221666 239982 223338 240038
rect 223506 239982 225178 240038
rect 225346 239982 227018 240038
rect 227186 239982 228858 240038
rect 229026 239982 230698 240038
rect 230866 239982 232538 240038
rect 232706 239982 234378 240038
rect 234546 239982 236218 240038
rect 236386 239982 237874 240038
rect 572 856 237986 239982
rect 682 800 2170 856
rect 2338 800 4010 856
rect 4178 800 5850 856
rect 6018 800 7690 856
rect 7858 800 9530 856
rect 9698 800 11370 856
rect 11538 800 13210 856
rect 13378 800 15050 856
rect 15218 800 16890 856
rect 17058 800 18730 856
rect 18898 800 20570 856
rect 20738 800 22410 856
rect 22578 800 24250 856
rect 24418 800 26090 856
rect 26258 800 27930 856
rect 28098 800 29770 856
rect 29938 800 31610 856
rect 31778 800 33450 856
rect 33618 800 35290 856
rect 35458 800 37130 856
rect 37298 800 38970 856
rect 39138 800 40626 856
rect 40794 800 42466 856
rect 42634 800 44306 856
rect 44474 800 46146 856
rect 46314 800 47986 856
rect 48154 800 49826 856
rect 49994 800 51666 856
rect 51834 800 53506 856
rect 53674 800 55346 856
rect 55514 800 57186 856
rect 57354 800 59026 856
rect 59194 800 60866 856
rect 61034 800 62706 856
rect 62874 800 64546 856
rect 64714 800 66386 856
rect 66554 800 68226 856
rect 68394 800 70066 856
rect 70234 800 71906 856
rect 72074 800 73746 856
rect 73914 800 75586 856
rect 75754 800 77426 856
rect 77594 800 79266 856
rect 79434 800 80922 856
rect 81090 800 82762 856
rect 82930 800 84602 856
rect 84770 800 86442 856
rect 86610 800 88282 856
rect 88450 800 90122 856
rect 90290 800 91962 856
rect 92130 800 93802 856
rect 93970 800 95642 856
rect 95810 800 97482 856
rect 97650 800 99322 856
rect 99490 800 101162 856
rect 101330 800 103002 856
rect 103170 800 104842 856
rect 105010 800 106682 856
rect 106850 800 108522 856
rect 108690 800 110362 856
rect 110530 800 112202 856
rect 112370 800 114042 856
rect 114210 800 115882 856
rect 116050 800 117722 856
rect 117890 800 119562 856
rect 119730 800 121218 856
rect 121386 800 123058 856
rect 123226 800 124898 856
rect 125066 800 126738 856
rect 126906 800 128578 856
rect 128746 800 130418 856
rect 130586 800 132258 856
rect 132426 800 134098 856
rect 134266 800 135938 856
rect 136106 800 137778 856
rect 137946 800 139618 856
rect 139786 800 141458 856
rect 141626 800 143298 856
rect 143466 800 145138 856
rect 145306 800 146978 856
rect 147146 800 148818 856
rect 148986 800 150658 856
rect 150826 800 152498 856
rect 152666 800 154338 856
rect 154506 800 156178 856
rect 156346 800 158018 856
rect 158186 800 159858 856
rect 160026 800 161514 856
rect 161682 800 163354 856
rect 163522 800 165194 856
rect 165362 800 167034 856
rect 167202 800 168874 856
rect 169042 800 170714 856
rect 170882 800 172554 856
rect 172722 800 174394 856
rect 174562 800 176234 856
rect 176402 800 178074 856
rect 178242 800 179914 856
rect 180082 800 181754 856
rect 181922 800 183594 856
rect 183762 800 185434 856
rect 185602 800 187274 856
rect 187442 800 189114 856
rect 189282 800 190954 856
rect 191122 800 192794 856
rect 192962 800 194634 856
rect 194802 800 196474 856
rect 196642 800 198314 856
rect 198482 800 200154 856
rect 200322 800 201810 856
rect 201978 800 203650 856
rect 203818 800 205490 856
rect 205658 800 207330 856
rect 207498 800 209170 856
rect 209338 800 211010 856
rect 211178 800 212850 856
rect 213018 800 214690 856
rect 214858 800 216530 856
rect 216698 800 218370 856
rect 218538 800 220210 856
rect 220378 800 222050 856
rect 222218 800 223890 856
rect 224058 800 225730 856
rect 225898 800 227570 856
rect 227738 800 229410 856
rect 229578 800 231250 856
rect 231418 800 233090 856
rect 233258 800 234930 856
rect 235098 800 236770 856
rect 236938 800 237986 856
<< metal3 >>
rect 0 238824 800 238944
rect 237894 237192 238694 237312
rect 0 236376 800 236496
rect 237894 234472 238694 234592
rect 0 233656 800 233776
rect 237894 231752 238694 231872
rect 0 230936 800 231056
rect 237894 229032 238694 229152
rect 0 228216 800 228336
rect 237894 226312 238694 226432
rect 0 225496 800 225616
rect 237894 223592 238694 223712
rect 0 222776 800 222896
rect 237894 220872 238694 220992
rect 0 220056 800 220176
rect 237894 218152 238694 218272
rect 0 217336 800 217456
rect 237894 215432 238694 215552
rect 0 214616 800 214736
rect 237894 212712 238694 212832
rect 0 211896 800 212016
rect 237894 209992 238694 210112
rect 0 209176 800 209296
rect 237894 207272 238694 207392
rect 0 206456 800 206576
rect 237894 204552 238694 204672
rect 0 203736 800 203856
rect 237894 201832 238694 201952
rect 0 201016 800 201136
rect 237894 199112 238694 199232
rect 0 198296 800 198416
rect 237894 196392 238694 196512
rect 0 195576 800 195696
rect 237894 193672 238694 193792
rect 0 192856 800 192976
rect 237894 190952 238694 191072
rect 0 190136 800 190256
rect 237894 188232 238694 188352
rect 0 187416 800 187536
rect 237894 185512 238694 185632
rect 0 184696 800 184816
rect 237894 182792 238694 182912
rect 0 181976 800 182096
rect 237894 180344 238694 180464
rect 0 179256 800 179376
rect 237894 177624 238694 177744
rect 0 176808 800 176928
rect 237894 174904 238694 175024
rect 0 174088 800 174208
rect 237894 172184 238694 172304
rect 0 171368 800 171488
rect 237894 169464 238694 169584
rect 0 168648 800 168768
rect 237894 166744 238694 166864
rect 0 165928 800 166048
rect 237894 164024 238694 164144
rect 0 163208 800 163328
rect 237894 161304 238694 161424
rect 0 160488 800 160608
rect 237894 158584 238694 158704
rect 0 157768 800 157888
rect 237894 155864 238694 155984
rect 0 155048 800 155168
rect 237894 153144 238694 153264
rect 0 152328 800 152448
rect 237894 150424 238694 150544
rect 0 149608 800 149728
rect 237894 147704 238694 147824
rect 0 146888 800 147008
rect 237894 144984 238694 145104
rect 0 144168 800 144288
rect 237894 142264 238694 142384
rect 0 141448 800 141568
rect 237894 139544 238694 139664
rect 0 138728 800 138848
rect 237894 136824 238694 136944
rect 0 136008 800 136128
rect 237894 134104 238694 134224
rect 0 133288 800 133408
rect 237894 131384 238694 131504
rect 0 130568 800 130688
rect 237894 128664 238694 128784
rect 0 127848 800 127968
rect 237894 125944 238694 126064
rect 0 125128 800 125248
rect 237894 123224 238694 123344
rect 0 122408 800 122528
rect 237894 120776 238694 120896
rect 0 119688 800 119808
rect 237894 118056 238694 118176
rect 0 117240 800 117360
rect 237894 115336 238694 115456
rect 0 114520 800 114640
rect 237894 112616 238694 112736
rect 0 111800 800 111920
rect 237894 109896 238694 110016
rect 0 109080 800 109200
rect 237894 107176 238694 107296
rect 0 106360 800 106480
rect 237894 104456 238694 104576
rect 0 103640 800 103760
rect 237894 101736 238694 101856
rect 0 100920 800 101040
rect 237894 99016 238694 99136
rect 0 98200 800 98320
rect 237894 96296 238694 96416
rect 0 95480 800 95600
rect 237894 93576 238694 93696
rect 0 92760 800 92880
rect 237894 90856 238694 90976
rect 0 90040 800 90160
rect 237894 88136 238694 88256
rect 0 87320 800 87440
rect 237894 85416 238694 85536
rect 0 84600 800 84720
rect 237894 82696 238694 82816
rect 0 81880 800 82000
rect 237894 79976 238694 80096
rect 0 79160 800 79280
rect 237894 77256 238694 77376
rect 0 76440 800 76560
rect 237894 74536 238694 74656
rect 0 73720 800 73840
rect 237894 71816 238694 71936
rect 0 71000 800 71120
rect 237894 69096 238694 69216
rect 0 68280 800 68400
rect 237894 66376 238694 66496
rect 0 65560 800 65680
rect 237894 63656 238694 63776
rect 0 62840 800 62960
rect 237894 61208 238694 61328
rect 0 60120 800 60240
rect 237894 58488 238694 58608
rect 0 57672 800 57792
rect 237894 55768 238694 55888
rect 0 54952 800 55072
rect 237894 53048 238694 53168
rect 0 52232 800 52352
rect 237894 50328 238694 50448
rect 0 49512 800 49632
rect 237894 47608 238694 47728
rect 0 46792 800 46912
rect 237894 44888 238694 45008
rect 0 44072 800 44192
rect 237894 42168 238694 42288
rect 0 41352 800 41472
rect 237894 39448 238694 39568
rect 0 38632 800 38752
rect 237894 36728 238694 36848
rect 0 35912 800 36032
rect 237894 34008 238694 34128
rect 0 33192 800 33312
rect 237894 31288 238694 31408
rect 0 30472 800 30592
rect 237894 28568 238694 28688
rect 0 27752 800 27872
rect 237894 25848 238694 25968
rect 0 25032 800 25152
rect 237894 23128 238694 23248
rect 0 22312 800 22432
rect 237894 20408 238694 20528
rect 0 19592 800 19712
rect 237894 17688 238694 17808
rect 0 16872 800 16992
rect 237894 14968 238694 15088
rect 0 14152 800 14272
rect 237894 12248 238694 12368
rect 0 11432 800 11552
rect 237894 9528 238694 9648
rect 0 8712 800 8832
rect 237894 6808 238694 6928
rect 0 5992 800 6112
rect 237894 4088 238694 4208
rect 0 3272 800 3392
rect 237894 1640 238694 1760
<< obsm3 >>
rect 880 238744 237991 238917
rect 798 237392 237991 238744
rect 798 237112 237814 237392
rect 798 236576 237991 237112
rect 880 236296 237991 236576
rect 798 234672 237991 236296
rect 798 234392 237814 234672
rect 798 233856 237991 234392
rect 880 233576 237991 233856
rect 798 231952 237991 233576
rect 798 231672 237814 231952
rect 798 231136 237991 231672
rect 880 230856 237991 231136
rect 798 229232 237991 230856
rect 798 228952 237814 229232
rect 798 228416 237991 228952
rect 880 228136 237991 228416
rect 798 226512 237991 228136
rect 798 226232 237814 226512
rect 798 225696 237991 226232
rect 880 225416 237991 225696
rect 798 223792 237991 225416
rect 798 223512 237814 223792
rect 798 222976 237991 223512
rect 880 222696 237991 222976
rect 798 221072 237991 222696
rect 798 220792 237814 221072
rect 798 220256 237991 220792
rect 880 219976 237991 220256
rect 798 218352 237991 219976
rect 798 218072 237814 218352
rect 798 217536 237991 218072
rect 880 217256 237991 217536
rect 798 215632 237991 217256
rect 798 215352 237814 215632
rect 798 214816 237991 215352
rect 880 214536 237991 214816
rect 798 212912 237991 214536
rect 798 212632 237814 212912
rect 798 212096 237991 212632
rect 880 211816 237991 212096
rect 798 210192 237991 211816
rect 798 209912 237814 210192
rect 798 209376 237991 209912
rect 880 209096 237991 209376
rect 798 207472 237991 209096
rect 798 207192 237814 207472
rect 798 206656 237991 207192
rect 880 206376 237991 206656
rect 798 204752 237991 206376
rect 798 204472 237814 204752
rect 798 203936 237991 204472
rect 880 203656 237991 203936
rect 798 202032 237991 203656
rect 798 201752 237814 202032
rect 798 201216 237991 201752
rect 880 200936 237991 201216
rect 798 199312 237991 200936
rect 798 199032 237814 199312
rect 798 198496 237991 199032
rect 880 198216 237991 198496
rect 798 196592 237991 198216
rect 798 196312 237814 196592
rect 798 195776 237991 196312
rect 880 195496 237991 195776
rect 798 193872 237991 195496
rect 798 193592 237814 193872
rect 798 193056 237991 193592
rect 880 192776 237991 193056
rect 798 191152 237991 192776
rect 798 190872 237814 191152
rect 798 190336 237991 190872
rect 880 190056 237991 190336
rect 798 188432 237991 190056
rect 798 188152 237814 188432
rect 798 187616 237991 188152
rect 880 187336 237991 187616
rect 798 185712 237991 187336
rect 798 185432 237814 185712
rect 798 184896 237991 185432
rect 880 184616 237991 184896
rect 798 182992 237991 184616
rect 798 182712 237814 182992
rect 798 182176 237991 182712
rect 880 181896 237991 182176
rect 798 180544 237991 181896
rect 798 180264 237814 180544
rect 798 179456 237991 180264
rect 880 179176 237991 179456
rect 798 177824 237991 179176
rect 798 177544 237814 177824
rect 798 177008 237991 177544
rect 880 176728 237991 177008
rect 798 175104 237991 176728
rect 798 174824 237814 175104
rect 798 174288 237991 174824
rect 880 174008 237991 174288
rect 798 172384 237991 174008
rect 798 172104 237814 172384
rect 798 171568 237991 172104
rect 880 171288 237991 171568
rect 798 169664 237991 171288
rect 798 169384 237814 169664
rect 798 168848 237991 169384
rect 880 168568 237991 168848
rect 798 166944 237991 168568
rect 798 166664 237814 166944
rect 798 166128 237991 166664
rect 880 165848 237991 166128
rect 798 164224 237991 165848
rect 798 163944 237814 164224
rect 798 163408 237991 163944
rect 880 163128 237991 163408
rect 798 161504 237991 163128
rect 798 161224 237814 161504
rect 798 160688 237991 161224
rect 880 160408 237991 160688
rect 798 158784 237991 160408
rect 798 158504 237814 158784
rect 798 157968 237991 158504
rect 880 157688 237991 157968
rect 798 156064 237991 157688
rect 798 155784 237814 156064
rect 798 155248 237991 155784
rect 880 154968 237991 155248
rect 798 153344 237991 154968
rect 798 153064 237814 153344
rect 798 152528 237991 153064
rect 880 152248 237991 152528
rect 798 150624 237991 152248
rect 798 150344 237814 150624
rect 798 149808 237991 150344
rect 880 149528 237991 149808
rect 798 147904 237991 149528
rect 798 147624 237814 147904
rect 798 147088 237991 147624
rect 880 146808 237991 147088
rect 798 145184 237991 146808
rect 798 144904 237814 145184
rect 798 144368 237991 144904
rect 880 144088 237991 144368
rect 798 142464 237991 144088
rect 798 142184 237814 142464
rect 798 141648 237991 142184
rect 880 141368 237991 141648
rect 798 139744 237991 141368
rect 798 139464 237814 139744
rect 798 138928 237991 139464
rect 880 138648 237991 138928
rect 798 137024 237991 138648
rect 798 136744 237814 137024
rect 798 136208 237991 136744
rect 880 135928 237991 136208
rect 798 134304 237991 135928
rect 798 134024 237814 134304
rect 798 133488 237991 134024
rect 880 133208 237991 133488
rect 798 131584 237991 133208
rect 798 131304 237814 131584
rect 798 130768 237991 131304
rect 880 130488 237991 130768
rect 798 128864 237991 130488
rect 798 128584 237814 128864
rect 798 128048 237991 128584
rect 880 127768 237991 128048
rect 798 126144 237991 127768
rect 798 125864 237814 126144
rect 798 125328 237991 125864
rect 880 125048 237991 125328
rect 798 123424 237991 125048
rect 798 123144 237814 123424
rect 798 122608 237991 123144
rect 880 122328 237991 122608
rect 798 120976 237991 122328
rect 798 120696 237814 120976
rect 798 119888 237991 120696
rect 880 119608 237991 119888
rect 798 118256 237991 119608
rect 798 117976 237814 118256
rect 798 117440 237991 117976
rect 880 117160 237991 117440
rect 798 115536 237991 117160
rect 798 115256 237814 115536
rect 798 114720 237991 115256
rect 880 114440 237991 114720
rect 798 112816 237991 114440
rect 798 112536 237814 112816
rect 798 112000 237991 112536
rect 880 111720 237991 112000
rect 798 110096 237991 111720
rect 798 109816 237814 110096
rect 798 109280 237991 109816
rect 880 109000 237991 109280
rect 798 107376 237991 109000
rect 798 107096 237814 107376
rect 798 106560 237991 107096
rect 880 106280 237991 106560
rect 798 104656 237991 106280
rect 798 104376 237814 104656
rect 798 103840 237991 104376
rect 880 103560 237991 103840
rect 798 101936 237991 103560
rect 798 101656 237814 101936
rect 798 101120 237991 101656
rect 880 100840 237991 101120
rect 798 99216 237991 100840
rect 798 98936 237814 99216
rect 798 98400 237991 98936
rect 880 98120 237991 98400
rect 798 96496 237991 98120
rect 798 96216 237814 96496
rect 798 95680 237991 96216
rect 880 95400 237991 95680
rect 798 93776 237991 95400
rect 798 93496 237814 93776
rect 798 92960 237991 93496
rect 880 92680 237991 92960
rect 798 91056 237991 92680
rect 798 90776 237814 91056
rect 798 90240 237991 90776
rect 880 89960 237991 90240
rect 798 88336 237991 89960
rect 798 88056 237814 88336
rect 798 87520 237991 88056
rect 880 87240 237991 87520
rect 798 85616 237991 87240
rect 798 85336 237814 85616
rect 798 84800 237991 85336
rect 880 84520 237991 84800
rect 798 82896 237991 84520
rect 798 82616 237814 82896
rect 798 82080 237991 82616
rect 880 81800 237991 82080
rect 798 80176 237991 81800
rect 798 79896 237814 80176
rect 798 79360 237991 79896
rect 880 79080 237991 79360
rect 798 77456 237991 79080
rect 798 77176 237814 77456
rect 798 76640 237991 77176
rect 880 76360 237991 76640
rect 798 74736 237991 76360
rect 798 74456 237814 74736
rect 798 73920 237991 74456
rect 880 73640 237991 73920
rect 798 72016 237991 73640
rect 798 71736 237814 72016
rect 798 71200 237991 71736
rect 880 70920 237991 71200
rect 798 69296 237991 70920
rect 798 69016 237814 69296
rect 798 68480 237991 69016
rect 880 68200 237991 68480
rect 798 66576 237991 68200
rect 798 66296 237814 66576
rect 798 65760 237991 66296
rect 880 65480 237991 65760
rect 798 63856 237991 65480
rect 798 63576 237814 63856
rect 798 63040 237991 63576
rect 880 62760 237991 63040
rect 798 61408 237991 62760
rect 798 61128 237814 61408
rect 798 60320 237991 61128
rect 880 60040 237991 60320
rect 798 58688 237991 60040
rect 798 58408 237814 58688
rect 798 57872 237991 58408
rect 880 57592 237991 57872
rect 798 55968 237991 57592
rect 798 55688 237814 55968
rect 798 55152 237991 55688
rect 880 54872 237991 55152
rect 798 53248 237991 54872
rect 798 52968 237814 53248
rect 798 52432 237991 52968
rect 880 52152 237991 52432
rect 798 50528 237991 52152
rect 798 50248 237814 50528
rect 798 49712 237991 50248
rect 880 49432 237991 49712
rect 798 47808 237991 49432
rect 798 47528 237814 47808
rect 798 46992 237991 47528
rect 880 46712 237991 46992
rect 798 45088 237991 46712
rect 798 44808 237814 45088
rect 798 44272 237991 44808
rect 880 43992 237991 44272
rect 798 42368 237991 43992
rect 798 42088 237814 42368
rect 798 41552 237991 42088
rect 880 41272 237991 41552
rect 798 39648 237991 41272
rect 798 39368 237814 39648
rect 798 38832 237991 39368
rect 880 38552 237991 38832
rect 798 36928 237991 38552
rect 798 36648 237814 36928
rect 798 36112 237991 36648
rect 880 35832 237991 36112
rect 798 34208 237991 35832
rect 798 33928 237814 34208
rect 798 33392 237991 33928
rect 880 33112 237991 33392
rect 798 31488 237991 33112
rect 798 31208 237814 31488
rect 798 30672 237991 31208
rect 880 30392 237991 30672
rect 798 28768 237991 30392
rect 798 28488 237814 28768
rect 798 27952 237991 28488
rect 880 27672 237991 27952
rect 798 26048 237991 27672
rect 798 25768 237814 26048
rect 798 25232 237991 25768
rect 880 24952 237991 25232
rect 798 23328 237991 24952
rect 798 23048 237814 23328
rect 798 22512 237991 23048
rect 880 22232 237991 22512
rect 798 20608 237991 22232
rect 798 20328 237814 20608
rect 798 19792 237991 20328
rect 880 19512 237991 19792
rect 798 17888 237991 19512
rect 798 17608 237814 17888
rect 798 17072 237991 17608
rect 880 16792 237991 17072
rect 798 15168 237991 16792
rect 798 14888 237814 15168
rect 798 14352 237991 14888
rect 880 14072 237991 14352
rect 798 12448 237991 14072
rect 798 12168 237814 12448
rect 798 11632 237991 12168
rect 880 11352 237991 11632
rect 798 9728 237991 11352
rect 798 9448 237814 9728
rect 798 8912 237991 9448
rect 880 8632 237991 8912
rect 798 7008 237991 8632
rect 798 6728 237814 7008
rect 798 6192 237991 6728
rect 880 5912 237991 6192
rect 798 4288 237991 5912
rect 798 4008 237814 4288
rect 798 3472 237991 4008
rect 880 3192 237991 3472
rect 798 1840 237991 3192
rect 798 1667 237814 1840
<< metal4 >>
rect 4208 2128 4528 238320
rect 19568 2128 19888 238320
<< obsm4 >>
rect 2635 2128 4128 238320
rect 4608 2128 19488 238320
rect 19968 2128 234928 238320
<< labels >>
rlabel metal2 s 34794 240038 34850 240838 6 clk
port 1 nsew default input
rlabel metal2 s 225234 240038 225290 240838 6 d_in[0]
port 2 nsew default input
rlabel metal2 s 7194 240038 7250 240838 6 d_in[10]
port 3 nsew default input
rlabel metal3 s 237894 9528 238694 9648 6 d_in[11]
port 4 nsew default input
rlabel metal2 s 172610 0 172666 800 6 d_in[12]
port 5 nsew default input
rlabel metal3 s 0 49512 800 49632 6 d_in[13]
port 6 nsew default input
rlabel metal2 s 230754 240038 230810 240838 6 d_in[14]
port 7 nsew default input
rlabel metal2 s 66442 0 66498 800 6 d_in[15]
port 8 nsew default input
rlabel metal3 s 0 163208 800 163328 6 d_in[16]
port 9 nsew default input
rlabel metal3 s 237894 79976 238694 80096 6 d_in[17]
port 10 nsew default input
rlabel metal3 s 0 87320 800 87440 6 d_in[18]
port 11 nsew default input
rlabel metal3 s 237894 204552 238694 204672 6 d_in[19]
port 12 nsew default input
rlabel metal2 s 22466 0 22522 800 6 d_in[1]
port 13 nsew default input
rlabel metal2 s 164698 240038 164754 240838 6 d_in[20]
port 14 nsew default input
rlabel metal2 s 60922 0 60978 800 6 d_in[21]
port 15 nsew default input
rlabel metal2 s 1674 240038 1730 240838 6 d_in[22]
port 16 nsew default input
rlabel metal3 s 237894 118056 238694 118176 6 d_in[23]
port 17 nsew default input
rlabel metal2 s 86498 0 86554 800 6 d_in[2]
port 18 nsew default input
rlabel metal2 s 35346 0 35402 800 6 d_in[3]
port 19 nsew default input
rlabel metal3 s 0 146888 800 147008 6 d_in[4]
port 20 nsew default input
rlabel metal2 s 131762 240038 131818 240838 6 d_in[5]
port 21 nsew default input
rlabel metal2 s 71962 0 72018 800 6 d_in[6]
port 22 nsew default input
rlabel metal2 s 71410 240038 71466 240838 6 d_in[7]
port 23 nsew default input
rlabel metal3 s 237894 71816 238694 71936 6 d_in[8]
port 24 nsew default input
rlabel metal3 s 0 84600 800 84720 6 d_in[9]
port 25 nsew default input
rlabel metal3 s 0 60120 800 60240 6 d_out[0]
port 26 nsew default output
rlabel metal3 s 0 106360 800 106480 6 d_out[100]
port 27 nsew default output
rlabel metal3 s 0 73720 800 73840 6 d_out[101]
port 28 nsew default output
rlabel metal2 s 150714 0 150770 800 6 d_out[102]
port 29 nsew default output
rlabel metal2 s 126242 240038 126298 240838 6 d_out[103]
port 30 nsew default output
rlabel metal2 s 67730 240038 67786 240838 6 d_out[104]
port 31 nsew default output
rlabel metal2 s 183098 240038 183154 240838 6 d_out[105]
port 32 nsew default output
rlabel metal2 s 121274 0 121330 800 6 d_out[106]
port 33 nsew default output
rlabel metal2 s 48042 0 48098 800 6 d_out[107]
port 34 nsew default output
rlabel metal2 s 84106 240038 84162 240838 6 d_out[108]
port 35 nsew default output
rlabel metal3 s 0 155048 800 155168 6 d_out[109]
port 36 nsew default output
rlabel metal2 s 231306 0 231362 800 6 d_out[10]
port 37 nsew default output
rlabel metal3 s 237894 237192 238694 237312 6 d_out[110]
port 38 nsew default output
rlabel metal2 s 184938 240038 184994 240838 6 d_out[111]
port 39 nsew default output
rlabel metal2 s 106186 240038 106242 240838 6 d_out[112]
port 40 nsew default output
rlabel metal2 s 210514 240038 210570 240838 6 d_out[113]
port 41 nsew default output
rlabel metal3 s 0 90040 800 90160 6 d_out[114]
port 42 nsew default output
rlabel metal2 s 29274 240038 29330 240838 6 d_out[115]
port 43 nsew default output
rlabel metal2 s 59082 0 59138 800 6 d_out[116]
port 44 nsew default output
rlabel metal3 s 237894 158584 238694 158704 6 d_out[117]
port 45 nsew default output
rlabel metal2 s 75090 240038 75146 240838 6 d_out[118]
port 46 nsew default output
rlabel metal2 s 214194 240038 214250 240838 6 d_out[119]
port 47 nsew default output
rlabel metal2 s 236826 0 236882 800 6 d_out[11]
port 48 nsew default output
rlabel metal2 s 44362 0 44418 800 6 d_out[120]
port 49 nsew default output
rlabel metal3 s 0 16872 800 16992 6 d_out[121]
port 50 nsew default output
rlabel metal2 s 109866 240038 109922 240838 6 d_out[122]
port 51 nsew default output
rlabel metal3 s 0 222776 800 222896 6 d_out[123]
port 52 nsew default output
rlabel metal2 s 216034 240038 216090 240838 6 d_out[124]
port 53 nsew default output
rlabel metal3 s 0 149608 800 149728 6 d_out[125]
port 54 nsew default output
rlabel metal2 s 75642 0 75698 800 6 d_out[126]
port 55 nsew default output
rlabel metal3 s 237894 12248 238694 12368 6 d_out[127]
port 56 nsew default output
rlabel metal2 s 196530 0 196586 800 6 d_out[128]
port 57 nsew default output
rlabel metal2 s 80426 240038 80482 240838 6 d_out[129]
port 58 nsew default output
rlabel metal2 s 47490 240038 47546 240838 6 d_out[12]
port 59 nsew default output
rlabel metal3 s 237894 85416 238694 85536 6 d_out[130]
port 60 nsew default output
rlabel metal3 s 0 144168 800 144288 6 d_out[131]
port 61 nsew default output
rlabel metal2 s 168378 240038 168434 240838 6 d_out[132]
port 62 nsew default output
rlabel metal2 s 178130 0 178186 800 6 d_out[133]
port 63 nsew default output
rlabel metal2 s 203706 0 203762 800 6 d_out[134]
port 64 nsew default output
rlabel metal3 s 237894 220872 238694 220992 6 d_out[135]
port 65 nsew default output
rlabel metal2 s 49882 0 49938 800 6 d_out[136]
port 66 nsew default output
rlabel metal2 s 174450 0 174506 800 6 d_out[137]
port 67 nsew default output
rlabel metal2 s 95698 0 95754 800 6 d_out[138]
port 68 nsew default output
rlabel metal2 s 175738 240038 175794 240838 6 d_out[139]
port 69 nsew default output
rlabel metal2 s 111706 240038 111762 240838 6 d_out[13]
port 70 nsew default output
rlabel metal2 s 62210 240038 62266 240838 6 d_out[140]
port 71 nsew default output
rlabel metal3 s 0 33192 800 33312 6 d_out[141]
port 72 nsew default output
rlabel metal2 s 76930 240038 76986 240838 6 d_out[142]
port 73 nsew default output
rlabel metal2 s 156234 0 156290 800 6 d_out[143]
port 74 nsew default output
rlabel metal2 s 18234 240038 18290 240838 6 d_out[144]
port 75 nsew default output
rlabel metal2 s 64602 0 64658 800 6 d_out[145]
port 76 nsew default output
rlabel metal3 s 0 5992 800 6112 6 d_out[146]
port 77 nsew default output
rlabel metal3 s 0 57672 800 57792 6 d_out[147]
port 78 nsew default output
rlabel metal2 s 80978 0 81034 800 6 d_out[148]
port 79 nsew default output
rlabel metal2 s 227626 0 227682 800 6 d_out[149]
port 80 nsew default output
rlabel metal3 s 237894 1640 238694 1760 6 d_out[14]
port 81 nsew default output
rlabel metal2 s 190458 240038 190514 240838 6 d_out[150]
port 82 nsew default output
rlabel metal2 s 100666 240038 100722 240838 6 d_out[151]
port 83 nsew default output
rlabel metal3 s 237894 128664 238694 128784 6 d_out[152]
port 84 nsew default output
rlabel metal2 s 4066 0 4122 800 6 d_out[153]
port 85 nsew default output
rlabel metal2 s 31666 0 31722 800 6 d_out[154]
port 86 nsew default output
rlabel metal3 s 0 174088 800 174208 6 d_out[155]
port 87 nsew default output
rlabel metal2 s 36634 240038 36690 240838 6 d_out[156]
port 88 nsew default output
rlabel metal2 s 183650 0 183706 800 6 d_out[157]
port 89 nsew default output
rlabel metal2 s 37186 0 37242 800 6 d_out[158]
port 90 nsew default output
rlabel metal2 s 77482 0 77538 800 6 d_out[159]
port 91 nsew default output
rlabel metal3 s 237894 42168 238694 42288 6 d_out[15]
port 92 nsew default output
rlabel metal2 s 170218 240038 170274 240838 6 d_out[160]
port 93 nsew default output
rlabel metal3 s 0 206456 800 206576 6 d_out[161]
port 94 nsew default output
rlabel metal2 s 62762 0 62818 800 6 d_out[162]
port 95 nsew default output
rlabel metal3 s 0 8712 800 8832 6 d_out[163]
port 96 nsew default output
rlabel metal2 s 70122 0 70178 800 6 d_out[164]
port 97 nsew default output
rlabel metal2 s 53010 240038 53066 240838 6 d_out[165]
port 98 nsew default output
rlabel metal2 s 91466 240038 91522 240838 6 d_out[166]
port 99 nsew default output
rlabel metal3 s 0 100920 800 101040 6 d_out[167]
port 100 nsew default output
rlabel metal3 s 237894 185512 238694 185632 6 d_out[168]
port 101 nsew default output
rlabel metal3 s 0 184696 800 184816 6 d_out[169]
port 102 nsew default output
rlabel metal3 s 0 81880 800 82000 6 d_out[16]
port 103 nsew default output
rlabel metal2 s 69570 240038 69626 240838 6 d_out[170]
port 104 nsew default output
rlabel metal3 s 237894 201832 238694 201952 6 d_out[171]
port 105 nsew default output
rlabel metal3 s 237894 39448 238694 39568 6 d_out[172]
port 106 nsew default output
rlabel metal2 s 95146 240038 95202 240838 6 d_out[173]
port 107 nsew default output
rlabel metal3 s 0 192856 800 192976 6 d_out[174]
port 108 nsew default output
rlabel metal2 s 234434 240038 234490 240838 6 d_out[175]
port 109 nsew default output
rlabel metal2 s 200210 0 200266 800 6 d_out[176]
port 110 nsew default output
rlabel metal2 s 25594 240038 25650 240838 6 d_out[177]
port 111 nsew default output
rlabel metal2 s 82818 0 82874 800 6 d_out[178]
port 112 nsew default output
rlabel metal2 s 181810 0 181866 800 6 d_out[179]
port 113 nsew default output
rlabel metal2 s 176290 0 176346 800 6 d_out[17]
port 114 nsew default output
rlabel metal2 s 158074 0 158130 800 6 d_out[180]
port 115 nsew default output
rlabel metal3 s 237894 177624 238694 177744 6 d_out[181]
port 116 nsew default output
rlabel metal3 s 237894 125944 238694 126064 6 d_out[182]
port 117 nsew default output
rlabel metal3 s 0 35912 800 36032 6 d_out[183]
port 118 nsew default output
rlabel metal2 s 41970 240038 42026 240838 6 d_out[184]
port 119 nsew default output
rlabel metal3 s 0 201016 800 201136 6 d_out[185]
port 120 nsew default output
rlabel metal3 s 237894 25848 238694 25968 6 d_out[186]
port 121 nsew default output
rlabel metal3 s 237894 107176 238694 107296 6 d_out[187]
port 122 nsew default output
rlabel metal3 s 237894 223592 238694 223712 6 d_out[188]
port 123 nsew default output
rlabel metal2 s 60370 240038 60426 240838 6 d_out[189]
port 124 nsew default output
rlabel metal2 s 132314 0 132370 800 6 d_out[18]
port 125 nsew default output
rlabel metal2 s 117778 0 117834 800 6 d_out[190]
port 126 nsew default output
rlabel metal2 s 5906 0 5962 800 6 d_out[191]
port 127 nsew default output
rlabel metal2 s 191010 0 191066 800 6 d_out[19]
port 128 nsew default output
rlabel metal3 s 237894 50328 238694 50448 6 d_out[1]
port 129 nsew default output
rlabel metal3 s 237894 77256 238694 77376 6 d_out[20]
port 130 nsew default output
rlabel metal3 s 0 41352 800 41472 6 d_out[21]
port 131 nsew default output
rlabel metal2 s 188618 240038 188674 240838 6 d_out[22]
port 132 nsew default output
rlabel metal2 s 51722 0 51778 800 6 d_out[23]
port 133 nsew default output
rlabel metal3 s 0 236376 800 236496 6 d_out[24]
port 134 nsew default output
rlabel metal2 s 209226 0 209282 800 6 d_out[25]
port 135 nsew default output
rlabel metal2 s 20626 0 20682 800 6 d_out[26]
port 136 nsew default output
rlabel metal3 s 237894 58488 238694 58608 6 d_out[27]
port 137 nsew default output
rlabel metal3 s 0 111800 800 111920 6 d_out[28]
port 138 nsew default output
rlabel metal2 s 113546 240038 113602 240838 6 d_out[29]
port 139 nsew default output
rlabel metal3 s 0 165928 800 166048 6 d_out[2]
port 140 nsew default output
rlabel metal2 s 219714 240038 219770 240838 6 d_out[30]
port 141 nsew default output
rlabel metal2 s 157522 240038 157578 240838 6 d_out[31]
port 142 nsew default output
rlabel metal3 s 237894 112616 238694 112736 6 d_out[32]
port 143 nsew default output
rlabel metal2 s 133602 240038 133658 240838 6 d_out[33]
port 144 nsew default output
rlabel metal2 s 137834 0 137890 800 6 d_out[34]
port 145 nsew default output
rlabel metal2 s 78586 240038 78642 240838 6 d_out[35]
port 146 nsew default output
rlabel metal2 s 84658 0 84714 800 6 d_out[36]
port 147 nsew default output
rlabel metal2 s 79322 0 79378 800 6 d_out[37]
port 148 nsew default output
rlabel metal3 s 0 71000 800 71120 6 d_out[38]
port 149 nsew default output
rlabel metal3 s 237894 153144 238694 153264 6 d_out[39]
port 150 nsew default output
rlabel metal2 s 24306 0 24362 800 6 d_out[3]
port 151 nsew default output
rlabel metal3 s 237894 150424 238694 150544 6 d_out[40]
port 152 nsew default output
rlabel metal3 s 237894 88136 238694 88256 6 d_out[41]
port 153 nsew default output
rlabel metal2 s 23754 240038 23810 240838 6 d_out[42]
port 154 nsew default output
rlabel metal3 s 237894 199112 238694 199232 6 d_out[43]
port 155 nsew default output
rlabel metal2 s 212906 0 212962 800 6 d_out[44]
port 156 nsew default output
rlabel metal2 s 27986 0 28042 800 6 d_out[45]
port 157 nsew default output
rlabel metal2 s 98826 240038 98882 240838 6 d_out[46]
port 158 nsew default output
rlabel metal2 s 195978 240038 196034 240838 6 d_out[47]
port 159 nsew default output
rlabel metal2 s 159178 240038 159234 240838 6 d_out[48]
port 160 nsew default output
rlabel metal3 s 0 46792 800 46912 6 d_out[49]
port 161 nsew default output
rlabel metal2 s 115938 0 115994 800 6 d_out[4]
port 162 nsew default output
rlabel metal3 s 237894 196392 238694 196512 6 d_out[50]
port 163 nsew default output
rlabel metal3 s 0 27752 800 27872 6 d_out[51]
port 164 nsew default output
rlabel metal3 s 0 127848 800 127968 6 d_out[52]
port 165 nsew default output
rlabel metal2 s 99378 0 99434 800 6 d_out[53]
port 166 nsew default output
rlabel metal2 s 93306 240038 93362 240838 6 d_out[54]
port 167 nsew default output
rlabel metal2 s 217874 240038 217930 240838 6 d_out[55]
port 168 nsew default output
rlabel metal2 s 112258 0 112314 800 6 d_out[56]
port 169 nsew default output
rlabel metal2 s 137282 240038 137338 240838 6 d_out[57]
port 170 nsew default output
rlabel metal3 s 0 214616 800 214736 6 d_out[58]
port 171 nsew default output
rlabel metal2 s 185490 0 185546 800 6 d_out[59]
port 172 nsew default output
rlabel metal3 s 237894 142264 238694 142384 6 d_out[5]
port 173 nsew default output
rlabel metal2 s 120722 240038 120778 240838 6 d_out[60]
port 174 nsew default output
rlabel metal2 s 148322 240038 148378 240838 6 d_out[61]
port 175 nsew default output
rlabel metal2 s 26146 0 26202 800 6 d_out[62]
port 176 nsew default output
rlabel metal3 s 0 79160 800 79280 6 d_out[63]
port 177 nsew default output
rlabel metal3 s 0 176808 800 176928 6 d_out[64]
port 178 nsew default output
rlabel metal2 s 12714 240038 12770 240838 6 d_out[65]
port 179 nsew default output
rlabel metal3 s 237894 166744 238694 166864 6 d_out[66]
port 180 nsew default output
rlabel metal3 s 237894 188232 238694 188352 6 d_out[67]
port 181 nsew default output
rlabel metal3 s 0 181976 800 182096 6 d_out[68]
port 182 nsew default output
rlabel metal3 s 237894 180344 238694 180464 6 d_out[69]
port 183 nsew default output
rlabel metal2 s 101218 0 101274 800 6 d_out[6]
port 184 nsew default output
rlabel metal3 s 237894 31288 238694 31408 6 d_out[70]
port 185 nsew default output
rlabel metal3 s 0 220056 800 220176 6 d_out[71]
port 186 nsew default output
rlabel metal2 s 570 0 626 800 6 d_out[72]
port 187 nsew default output
rlabel metal2 s 142802 240038 142858 240838 6 d_out[73]
port 188 nsew default output
rlabel metal2 s 39026 0 39082 800 6 d_out[74]
port 189 nsew default output
rlabel metal2 s 18786 0 18842 800 6 d_out[75]
port 190 nsew default output
rlabel metal2 s 199474 240038 199530 240838 6 d_out[76]
port 191 nsew default output
rlabel metal3 s 0 233656 800 233776 6 d_out[77]
port 192 nsew default output
rlabel metal2 s 64050 240038 64106 240838 6 d_out[78]
port 193 nsew default output
rlabel metal2 s 104346 240038 104402 240838 6 d_out[79]
port 194 nsew default output
rlabel metal2 s 96986 240038 97042 240838 6 d_out[7]
port 195 nsew default output
rlabel metal3 s 237894 61208 238694 61328 6 d_out[80]
port 196 nsew default output
rlabel metal3 s 237894 104456 238694 104576 6 d_out[81]
port 197 nsew default output
rlabel metal2 s 233146 0 233202 800 6 d_out[82]
port 198 nsew default output
rlabel metal3 s 237894 209992 238694 210112 6 d_out[83]
port 199 nsew default output
rlabel metal2 s 3514 240038 3570 240838 6 d_out[84]
port 200 nsew default output
rlabel metal3 s 237894 136824 238694 136944 6 d_out[85]
port 201 nsew default output
rlabel metal3 s 0 228216 800 228336 6 d_out[86]
port 202 nsew default output
rlabel metal3 s 0 230936 800 231056 6 d_out[87]
port 203 nsew default output
rlabel metal3 s 237894 20408 238694 20528 6 d_out[88]
port 204 nsew default output
rlabel metal2 s 207386 0 207442 800 6 d_out[89]
port 205 nsew default output
rlabel metal2 s 223394 240038 223450 240838 6 d_out[8]
port 206 nsew default output
rlabel metal3 s 0 117240 800 117360 6 d_out[90]
port 207 nsew default output
rlabel metal3 s 0 211896 800 212016 6 d_out[91]
port 208 nsew default output
rlabel metal2 s 87786 240038 87842 240838 6 d_out[92]
port 209 nsew default output
rlabel metal3 s 0 179256 800 179376 6 d_out[93]
port 210 nsew default output
rlabel metal3 s 237894 34008 238694 34128 6 d_out[94]
port 211 nsew default output
rlabel metal2 s 82266 240038 82322 240838 6 d_out[95]
port 212 nsew default output
rlabel metal3 s 0 25032 800 25152 6 d_out[96]
port 213 nsew default output
rlabel metal2 s 152554 0 152610 800 6 d_out[97]
port 214 nsew default output
rlabel metal2 s 124954 0 125010 800 6 d_out[98]
port 215 nsew default output
rlabel metal2 s 237930 240038 237986 240838 6 d_out[99]
port 216 nsew default output
rlabel metal3 s 237894 155864 238694 155984 6 d_out[9]
port 217 nsew default output
rlabel metal3 s 237894 55768 238694 55888 6 dbg_gpr_ack
port 218 nsew default output
rlabel metal3 s 237894 74536 238694 74656 6 dbg_gpr_addr[0]
port 219 nsew default input
rlabel metal2 s 177578 240038 177634 240838 6 dbg_gpr_addr[1]
port 220 nsew default input
rlabel metal3 s 237894 28568 238694 28688 6 dbg_gpr_addr[2]
port 221 nsew default input
rlabel metal3 s 237894 115336 238694 115456 6 dbg_gpr_addr[3]
port 222 nsew default input
rlabel metal2 s 102506 240038 102562 240838 6 dbg_gpr_addr[4]
port 223 nsew default input
rlabel metal3 s 0 103640 800 103760 6 dbg_gpr_addr[5]
port 224 nsew default input
rlabel metal2 s 15106 0 15162 800 6 dbg_gpr_addr[6]
port 225 nsew default input
rlabel metal2 s 187330 0 187386 800 6 dbg_gpr_data[0]
port 226 nsew default output
rlabel metal3 s 237894 47608 238694 47728 6 dbg_gpr_data[10]
port 227 nsew default output
rlabel metal3 s 0 65560 800 65680 6 dbg_gpr_data[11]
port 228 nsew default output
rlabel metal3 s 237894 23128 238694 23248 6 dbg_gpr_data[12]
port 229 nsew default output
rlabel metal3 s 0 3272 800 3392 6 dbg_gpr_data[13]
port 230 nsew default output
rlabel metal3 s 237894 99016 238694 99136 6 dbg_gpr_data[14]
port 231 nsew default output
rlabel metal3 s 0 62840 800 62960 6 dbg_gpr_data[15]
port 232 nsew default output
rlabel metal2 s 32954 240038 33010 240838 6 dbg_gpr_data[16]
port 233 nsew default output
rlabel metal3 s 237894 69096 238694 69216 6 dbg_gpr_data[17]
port 234 nsew default output
rlabel metal2 s 53562 0 53618 800 6 dbg_gpr_data[18]
port 235 nsew default output
rlabel metal2 s 128634 0 128690 800 6 dbg_gpr_data[19]
port 236 nsew default output
rlabel metal2 s 173898 240038 173954 240838 6 dbg_gpr_data[1]
port 237 nsew default output
rlabel metal3 s 237894 193672 238694 193792 6 dbg_gpr_data[20]
port 238 nsew default output
rlabel metal2 s 73802 0 73858 800 6 dbg_gpr_data[21]
port 239 nsew default output
rlabel metal2 s 223946 0 224002 800 6 dbg_gpr_data[22]
port 240 nsew default output
rlabel metal2 s 172058 240038 172114 240838 6 dbg_gpr_data[23]
port 241 nsew default output
rlabel metal2 s 57242 0 57298 800 6 dbg_gpr_data[24]
port 242 nsew default output
rlabel metal2 s 154394 0 154450 800 6 dbg_gpr_data[25]
port 243 nsew default output
rlabel metal3 s 237894 82696 238694 82816 6 dbg_gpr_data[26]
port 244 nsew default output
rlabel metal3 s 237894 131384 238694 131504 6 dbg_gpr_data[27]
port 245 nsew default output
rlabel metal2 s 40682 0 40738 800 6 dbg_gpr_data[28]
port 246 nsew default output
rlabel metal2 s 16946 0 17002 800 6 dbg_gpr_data[29]
port 247 nsew default output
rlabel metal2 s 204994 240038 205050 240838 6 dbg_gpr_data[2]
port 248 nsew default output
rlabel metal2 s 42522 0 42578 800 6 dbg_gpr_data[30]
port 249 nsew default output
rlabel metal2 s 103058 0 103114 800 6 dbg_gpr_data[31]
port 250 nsew default output
rlabel metal3 s 0 195576 800 195696 6 dbg_gpr_data[32]
port 251 nsew default output
rlabel metal2 s 218426 0 218482 800 6 dbg_gpr_data[33]
port 252 nsew default output
rlabel metal2 s 161570 0 161626 800 6 dbg_gpr_data[34]
port 253 nsew default output
rlabel metal2 s 54850 240038 54906 240838 6 dbg_gpr_data[35]
port 254 nsew default output
rlabel metal2 s 167090 0 167146 800 6 dbg_gpr_data[36]
port 255 nsew default output
rlabel metal2 s 162858 240038 162914 240838 6 dbg_gpr_data[37]
port 256 nsew default output
rlabel metal2 s 194690 0 194746 800 6 dbg_gpr_data[38]
port 257 nsew default output
rlabel metal2 s 93858 0 93914 800 6 dbg_gpr_data[39]
port 258 nsew default output
rlabel metal2 s 40130 240038 40186 240838 6 dbg_gpr_data[3]
port 259 nsew default output
rlabel metal2 s 89626 240038 89682 240838 6 dbg_gpr_data[40]
port 260 nsew default output
rlabel metal2 s 222106 0 222162 800 6 dbg_gpr_data[41]
port 261 nsew default output
rlabel metal2 s 236274 240038 236330 240838 6 dbg_gpr_data[42]
port 262 nsew default output
rlabel metal2 s 206834 240038 206890 240838 6 dbg_gpr_data[43]
port 263 nsew default output
rlabel metal2 s 118882 240038 118938 240838 6 dbg_gpr_data[44]
port 264 nsew default output
rlabel metal2 s 58530 240038 58586 240838 6 dbg_gpr_data[45]
port 265 nsew default output
rlabel metal3 s 0 68280 800 68400 6 dbg_gpr_data[46]
port 266 nsew default output
rlabel metal2 s 21914 240038 21970 240838 6 dbg_gpr_data[47]
port 267 nsew default output
rlabel metal2 s 31114 240038 31170 240838 6 dbg_gpr_data[48]
port 268 nsew default output
rlabel metal2 s 104898 0 104954 800 6 dbg_gpr_data[49]
port 269 nsew default output
rlabel metal3 s 0 209176 800 209296 6 dbg_gpr_data[4]
port 270 nsew default output
rlabel metal3 s 237894 190952 238694 191072 6 dbg_gpr_data[50]
port 271 nsew default output
rlabel metal2 s 159914 0 159970 800 6 dbg_gpr_data[51]
port 272 nsew default output
rlabel metal3 s 237894 53048 238694 53168 6 dbg_gpr_data[52]
port 273 nsew default output
rlabel metal2 s 29826 0 29882 800 6 dbg_gpr_data[53]
port 274 nsew default output
rlabel metal3 s 0 157768 800 157888 6 dbg_gpr_data[54]
port 275 nsew default output
rlabel metal3 s 0 198296 800 198416 6 dbg_gpr_data[55]
port 276 nsew default output
rlabel metal2 s 126794 0 126850 800 6 dbg_gpr_data[56]
port 277 nsew default output
rlabel metal3 s 237894 90856 238694 90976 6 dbg_gpr_data[57]
port 278 nsew default output
rlabel metal3 s 0 14152 800 14272 6 dbg_gpr_data[58]
port 279 nsew default output
rlabel metal2 s 234986 0 235042 800 6 dbg_gpr_data[59]
port 280 nsew default output
rlabel metal2 s 139122 240038 139178 240838 6 dbg_gpr_data[5]
port 281 nsew default output
rlabel metal3 s 0 122408 800 122528 6 dbg_gpr_data[60]
port 282 nsew default output
rlabel metal2 s 117226 240038 117282 240838 6 dbg_gpr_data[61]
port 283 nsew default output
rlabel metal3 s 0 19592 800 19712 6 dbg_gpr_data[62]
port 284 nsew default output
rlabel metal2 s 155682 240038 155738 240838 6 dbg_gpr_data[63]
port 285 nsew default output
rlabel metal3 s 237894 229032 238694 229152 6 dbg_gpr_data[6]
port 286 nsew default output
rlabel metal2 s 51170 240038 51226 240838 6 dbg_gpr_data[7]
port 287 nsew default output
rlabel metal2 s 108026 240038 108082 240838 6 dbg_gpr_data[8]
port 288 nsew default output
rlabel metal2 s 181258 240038 181314 240838 6 dbg_gpr_data[9]
port 289 nsew default output
rlabel metal3 s 237894 147704 238694 147824 6 dbg_gpr_req
port 290 nsew default input
rlabel metal2 s 227074 240038 227130 240838 6 log_out[0]
port 291 nsew default output
rlabel metal2 s 55402 0 55458 800 6 log_out[10]
port 292 nsew default output
rlabel metal2 s 228914 240038 228970 240838 6 log_out[11]
port 293 nsew default output
rlabel metal2 s 9034 240038 9090 240838 6 log_out[12]
port 294 nsew default output
rlabel metal2 s 192850 0 192906 800 6 log_out[13]
port 295 nsew default output
rlabel metal3 s 0 238824 800 238944 6 log_out[14]
port 296 nsew default output
rlabel metal3 s 237894 123224 238694 123344 6 log_out[15]
port 297 nsew default output
rlabel metal3 s 237894 207272 238694 207392 6 log_out[16]
port 298 nsew default output
rlabel metal3 s 237894 169464 238694 169584 6 log_out[17]
port 299 nsew default output
rlabel metal2 s 165250 0 165306 800 6 log_out[18]
port 300 nsew default output
rlabel metal2 s 152002 240038 152058 240838 6 log_out[19]
port 301 nsew default output
rlabel metal3 s 237894 14968 238694 15088 6 log_out[1]
port 302 nsew default output
rlabel metal3 s 0 171368 800 171488 6 log_out[20]
port 303 nsew default output
rlabel metal2 s 130474 0 130530 800 6 log_out[21]
port 304 nsew default output
rlabel metal2 s 10874 240038 10930 240838 6 log_out[22]
port 305 nsew default output
rlabel metal3 s 0 225496 800 225616 6 log_out[23]
port 306 nsew default output
rlabel metal2 s 179418 240038 179474 240838 6 log_out[24]
port 307 nsew default output
rlabel metal3 s 0 52232 800 52352 6 log_out[25]
port 308 nsew default output
rlabel metal2 s 106738 0 106794 800 6 log_out[26]
port 309 nsew default output
rlabel metal2 s 97538 0 97594 800 6 log_out[27]
port 310 nsew default output
rlabel metal3 s 0 125128 800 125248 6 log_out[28]
port 311 nsew default output
rlabel metal2 s 73250 240038 73306 240838 6 log_out[29]
port 312 nsew default output
rlabel metal2 s 198370 0 198426 800 6 log_out[2]
port 313 nsew default output
rlabel metal2 s 163410 0 163466 800 6 log_out[30]
port 314 nsew default output
rlabel metal3 s 0 22312 800 22432 6 log_out[31]
port 315 nsew default output
rlabel metal3 s 237894 161304 238694 161424 6 log_out[32]
port 316 nsew default output
rlabel metal2 s 14554 240038 14610 240838 6 log_out[33]
port 317 nsew default output
rlabel metal2 s 134154 0 134210 800 6 log_out[34]
port 318 nsew default output
rlabel metal2 s 122562 240038 122618 240838 6 log_out[35]
port 319 nsew default output
rlabel metal2 s 33506 0 33562 800 6 log_out[36]
port 320 nsew default output
rlabel metal2 s 27434 240038 27490 240838 6 log_out[37]
port 321 nsew default output
rlabel metal3 s 0 190136 800 190256 6 log_out[38]
port 322 nsew default output
rlabel metal3 s 237894 234472 238694 234592 6 log_out[39]
port 323 nsew default output
rlabel metal2 s 147034 0 147090 800 6 log_out[3]
port 324 nsew default output
rlabel metal2 s 179970 0 180026 800 6 log_out[40]
port 325 nsew default output
rlabel metal2 s 135442 240038 135498 240838 6 log_out[41]
port 326 nsew default output
rlabel metal3 s 237894 96296 238694 96416 6 log_out[42]
port 327 nsew default output
rlabel metal3 s 0 168648 800 168768 6 log_out[43]
port 328 nsew default output
rlabel metal2 s 201314 240038 201370 240838 6 log_out[44]
port 329 nsew default output
rlabel metal2 s 90178 0 90234 800 6 log_out[45]
port 330 nsew default output
rlabel metal2 s 5354 240038 5410 240838 6 log_out[46]
port 331 nsew default output
rlabel metal3 s 0 187416 800 187536 6 log_out[47]
port 332 nsew default output
rlabel metal2 s 214746 0 214802 800 6 log_out[48]
port 333 nsew default output
rlabel metal2 s 110418 0 110474 800 6 log_out[49]
port 334 nsew default output
rlabel metal2 s 220266 0 220322 800 6 log_out[4]
port 335 nsew default output
rlabel metal3 s 237894 17688 238694 17808 6 log_out[50]
port 336 nsew default output
rlabel metal3 s 0 114520 800 114640 6 log_out[51]
port 337 nsew default output
rlabel metal3 s 0 30472 800 30592 6 log_out[52]
port 338 nsew default output
rlabel metal2 s 197818 240038 197874 240838 6 log_out[53]
port 339 nsew default output
rlabel metal3 s 237894 63656 238694 63776 6 log_out[54]
port 340 nsew default output
rlabel metal3 s 237894 139544 238694 139664 6 log_out[55]
port 341 nsew default output
rlabel metal3 s 237894 93576 238694 93696 6 log_out[56]
port 342 nsew default output
rlabel metal3 s 0 44072 800 44192 6 log_out[57]
port 343 nsew default output
rlabel metal2 s 65890 240038 65946 240838 6 log_out[58]
port 344 nsew default output
rlabel metal2 s 135994 0 136050 800 6 log_out[59]
port 345 nsew default output
rlabel metal3 s 237894 36728 238694 36848 6 log_out[5]
port 346 nsew default output
rlabel metal2 s 13266 0 13322 800 6 log_out[60]
port 347 nsew default output
rlabel metal3 s 237894 212712 238694 212832 6 log_out[61]
port 348 nsew default output
rlabel metal2 s 88338 0 88394 800 6 log_out[62]
port 349 nsew default output
rlabel metal2 s 108578 0 108634 800 6 log_out[63]
port 350 nsew default output
rlabel metal2 s 201866 0 201922 800 6 log_out[64]
port 351 nsew default output
rlabel metal2 s 16394 240038 16450 240838 6 log_out[65]
port 352 nsew default output
rlabel metal3 s 237894 6808 238694 6928 6 log_out[66]
port 353 nsew default output
rlabel metal2 s 192298 240038 192354 240838 6 log_out[67]
port 354 nsew default output
rlabel metal2 s 205546 0 205602 800 6 log_out[68]
port 355 nsew default output
rlabel metal2 s 43810 240038 43866 240838 6 log_out[69]
port 356 nsew default output
rlabel metal2 s 229466 0 229522 800 6 log_out[6]
port 357 nsew default output
rlabel metal3 s 0 109080 800 109200 6 log_out[70]
port 358 nsew default output
rlabel metal3 s 0 76440 800 76560 6 log_out[71]
port 359 nsew default output
rlabel metal3 s 237894 226312 238694 226432 6 log_out[7]
port 360 nsew default output
rlabel metal3 s 237894 4088 238694 4208 6 log_out[8]
port 361 nsew default output
rlabel metal2 s 208674 240038 208730 240838 6 log_out[9]
port 362 nsew default output
rlabel metal3 s 0 54952 800 55072 6 sim_dump
port 363 nsew default input
rlabel metal2 s 212354 240038 212410 240838 6 sim_dump_done
port 364 nsew default output
rlabel metal3 s 237894 101736 238694 101856 6 w_in[0]
port 365 nsew default input
rlabel metal2 s 124402 240038 124458 240838 6 w_in[10]
port 366 nsew default input
rlabel metal2 s 9586 0 9642 800 6 w_in[11]
port 367 nsew default input
rlabel metal2 s 56690 240038 56746 240838 6 w_in[12]
port 368 nsew default input
rlabel metal2 s 45650 240038 45706 240838 6 w_in[13]
port 369 nsew default input
rlabel metal3 s 0 130568 800 130688 6 w_in[14]
port 370 nsew default input
rlabel metal3 s 0 138728 800 138848 6 w_in[15]
port 371 nsew default input
rlabel metal2 s 140962 240038 141018 240838 6 w_in[16]
port 372 nsew default input
rlabel metal3 s 0 119688 800 119808 6 w_in[17]
port 373 nsew default input
rlabel metal2 s 114098 0 114154 800 6 w_in[18]
port 374 nsew default input
rlabel metal2 s 123114 0 123170 800 6 w_in[19]
port 375 nsew default input
rlabel metal2 s 186778 240038 186834 240838 6 w_in[1]
port 376 nsew default input
rlabel metal2 s 221554 240038 221610 240838 6 w_in[20]
port 377 nsew default input
rlabel metal2 s 11426 0 11482 800 6 w_in[21]
port 378 nsew default input
rlabel metal2 s 141514 0 141570 800 6 w_in[22]
port 379 nsew default input
rlabel metal2 s 129922 240038 129978 240838 6 w_in[23]
port 380 nsew default input
rlabel metal3 s 0 95480 800 95600 6 w_in[24]
port 381 nsew default input
rlabel metal2 s 166538 240038 166594 240838 6 w_in[25]
port 382 nsew default input
rlabel metal3 s 0 98200 800 98320 6 w_in[26]
port 383 nsew default input
rlabel metal3 s 0 217336 800 217456 6 w_in[27]
port 384 nsew default input
rlabel metal2 s 216586 0 216642 800 6 w_in[28]
port 385 nsew default input
rlabel metal2 s 148874 0 148930 800 6 w_in[29]
port 386 nsew default input
rlabel metal2 s 68282 0 68338 800 6 w_in[2]
port 387 nsew default input
rlabel metal2 s 7746 0 7802 800 6 w_in[30]
port 388 nsew default input
rlabel metal3 s 0 38632 800 38752 6 w_in[31]
port 389 nsew default input
rlabel metal3 s 0 141448 800 141568 6 w_in[32]
port 390 nsew default input
rlabel metal3 s 237894 215432 238694 215552 6 w_in[33]
port 391 nsew default input
rlabel metal2 s 189170 0 189226 800 6 w_in[34]
port 392 nsew default input
rlabel metal3 s 0 11432 800 11552 6 w_in[35]
port 393 nsew default input
rlabel metal3 s 0 203736 800 203856 6 w_in[36]
port 394 nsew default input
rlabel metal2 s 211066 0 211122 800 6 w_in[37]
port 395 nsew default input
rlabel metal3 s 237894 144984 238694 145104 6 w_in[38]
port 396 nsew default input
rlabel metal3 s 0 136008 800 136128 6 w_in[39]
port 397 nsew default input
rlabel metal3 s 237894 109896 238694 110016 6 w_in[3]
port 398 nsew default input
rlabel metal2 s 85946 240038 86002 240838 6 w_in[40]
port 399 nsew default input
rlabel metal3 s 237894 172184 238694 172304 6 w_in[41]
port 400 nsew default input
rlabel metal2 s 46202 0 46258 800 6 w_in[42]
port 401 nsew default input
rlabel metal3 s 237894 174904 238694 175024 6 w_in[43]
port 402 nsew default input
rlabel metal2 s 20074 240038 20130 240838 6 w_in[44]
port 403 nsew default input
rlabel metal3 s 237894 44888 238694 45008 6 w_in[45]
port 404 nsew default input
rlabel metal3 s 237894 218152 238694 218272 6 w_in[46]
port 405 nsew default input
rlabel metal3 s 237894 231752 238694 231872 6 w_in[47]
port 406 nsew default input
rlabel metal2 s 144642 240038 144698 240838 6 w_in[48]
port 407 nsew default input
rlabel metal3 s 0 160488 800 160608 6 w_in[49]
port 408 nsew default input
rlabel metal2 s 203154 240038 203210 240838 6 w_in[4]
port 409 nsew default input
rlabel metal2 s 232594 240038 232650 240838 6 w_in[50]
port 410 nsew default input
rlabel metal2 s 143354 0 143410 800 6 w_in[51]
port 411 nsew default input
rlabel metal2 s 194138 240038 194194 240838 6 w_in[52]
port 412 nsew default input
rlabel metal3 s 0 152328 800 152448 6 w_in[53]
port 413 nsew default input
rlabel metal3 s 237894 182792 238694 182912 6 w_in[54]
port 414 nsew default input
rlabel metal2 s 49330 240038 49386 240838 6 w_in[55]
port 415 nsew default input
rlabel metal2 s 153842 240038 153898 240838 6 w_in[56]
port 416 nsew default input
rlabel metal2 s 139674 0 139730 800 6 w_in[57]
port 417 nsew default input
rlabel metal2 s 92018 0 92074 800 6 w_in[58]
port 418 nsew default input
rlabel metal3 s 237894 134104 238694 134224 6 w_in[59]
port 419 nsew default input
rlabel metal2 s 168930 0 168986 800 6 w_in[5]
port 420 nsew default input
rlabel metal3 s 237894 164024 238694 164144 6 w_in[60]
port 421 nsew default input
rlabel metal2 s 170770 0 170826 800 6 w_in[61]
port 422 nsew default input
rlabel metal2 s 225786 0 225842 800 6 w_in[62]
port 423 nsew default input
rlabel metal2 s 2226 0 2282 800 6 w_in[63]
port 424 nsew default input
rlabel metal3 s 237894 66376 238694 66496 6 w_in[64]
port 425 nsew default input
rlabel metal3 s 237894 120776 238694 120896 6 w_in[65]
port 426 nsew default input
rlabel metal3 s 0 133288 800 133408 6 w_in[66]
port 427 nsew default input
rlabel metal2 s 119618 0 119674 800 6 w_in[67]
port 428 nsew default input
rlabel metal2 s 161018 240038 161074 240838 6 w_in[68]
port 429 nsew default input
rlabel metal3 s 0 92760 800 92880 6 w_in[69]
port 430 nsew default input
rlabel metal2 s 145194 0 145250 800 6 w_in[6]
port 431 nsew default input
rlabel metal2 s 150162 240038 150218 240838 6 w_in[70]
port 432 nsew default input
rlabel metal2 s 115386 240038 115442 240838 6 w_in[71]
port 433 nsew default input
rlabel metal2 s 38290 240038 38346 240838 6 w_in[7]
port 434 nsew default input
rlabel metal2 s 146482 240038 146538 240838 6 w_in[8]
port 435 nsew default input
rlabel metal2 s 128082 240038 128138 240838 6 w_in[9]
port 436 nsew default input
rlabel metal4 s 4208 2128 4528 238320 6 VPWR
port 437 nsew power input
rlabel metal4 s 19568 2128 19888 238320 6 VGND
port 438 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 238694 240838
string LEFview TRUE
<< end >>
